-- Generator : SpinalHDL v1.6.1    git head : 3bf789d53b1b5a36974196e2d591342e15ddf28c
-- Component : Muraxy
-- Git hash  : 349993b23578fff6714024d38b53d5ccdafe11fd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;

package pkg_enum is
  type Axi4ToApb3BridgePhase is (SETUP,ACCESS_1,RESPONSE);
  type UartStopType is (ONE,TWO);
  type UartParityType is (NONE,EVEN,ODD);
  type UartCtrlTxState is (IDLE,START,DATA,PARITY,STOP);
  type UartCtrlRxState is (IDLE,START,DATA,PARITY,STOP);
  type EnvCtrlEnum is (NONE,XRET);
  type BranchCtrlEnum is (INC,B,JAL,JALR);
  type ShiftCtrlEnum is (DISABLE_1,SLL_1,SRL_1,SRA_1);
  type AluBitwiseCtrlEnum is (XOR_1,OR_1,AND_1);
  type Src2CtrlEnum is (RS,IMI,IMS,PC);
  type AluCtrlEnum is (ADD_SUB,SLT_SLTU,BITWISE);
  type Src1CtrlEnum is (RS,IMU,PC_INCREMENT,URS1);

  function pkg_mux (sel : std_logic; one : Axi4ToApb3BridgePhase; zero : Axi4ToApb3BridgePhase) return Axi4ToApb3BridgePhase;
  function pkg_toStdLogicVector_native (value : Axi4ToApb3BridgePhase) return std_logic_vector;
  function pkg_toAxi4ToApb3BridgePhase_native (value : std_logic_vector(1 downto 0)) return Axi4ToApb3BridgePhase;
  function pkg_mux (sel : std_logic; one : UartStopType; zero : UartStopType) return UartStopType;
  subtype UartStopType_seq_type is std_logic_vector(0 downto 0);
  constant UartStopType_seq_ONE : UartStopType_seq_type := "0";
  constant UartStopType_seq_TWO : UartStopType_seq_type := "1";

  function pkg_mux (sel : std_logic; one : UartParityType; zero : UartParityType) return UartParityType;
  subtype UartParityType_seq_type is std_logic_vector(1 downto 0);
  constant UartParityType_seq_NONE : UartParityType_seq_type := "00";
  constant UartParityType_seq_EVEN : UartParityType_seq_type := "01";
  constant UartParityType_seq_ODD : UartParityType_seq_type := "10";

  function pkg_mux (sel : std_logic; one : UartCtrlTxState; zero : UartCtrlTxState) return UartCtrlTxState;
  function pkg_toStdLogicVector_native (value : UartCtrlTxState) return std_logic_vector;
  function pkg_toUartCtrlTxState_native (value : std_logic_vector(2 downto 0)) return UartCtrlTxState;
  function pkg_mux (sel : std_logic; one : UartCtrlRxState; zero : UartCtrlRxState) return UartCtrlRxState;
  function pkg_toStdLogicVector_native (value : UartCtrlRxState) return std_logic_vector;
  function pkg_toUartCtrlRxState_native (value : std_logic_vector(2 downto 0)) return UartCtrlRxState;
  function pkg_mux (sel : std_logic; one : EnvCtrlEnum; zero : EnvCtrlEnum) return EnvCtrlEnum;
  subtype EnvCtrlEnum_seq_type is std_logic_vector(0 downto 0);
  constant EnvCtrlEnum_seq_NONE : EnvCtrlEnum_seq_type := "0";
  constant EnvCtrlEnum_seq_XRET : EnvCtrlEnum_seq_type := "1";

  function pkg_mux (sel : std_logic; one : BranchCtrlEnum; zero : BranchCtrlEnum) return BranchCtrlEnum;
  subtype BranchCtrlEnum_seq_type is std_logic_vector(1 downto 0);
  constant BranchCtrlEnum_seq_INC : BranchCtrlEnum_seq_type := "00";
  constant BranchCtrlEnum_seq_B : BranchCtrlEnum_seq_type := "01";
  constant BranchCtrlEnum_seq_JAL : BranchCtrlEnum_seq_type := "10";
  constant BranchCtrlEnum_seq_JALR : BranchCtrlEnum_seq_type := "11";

  function pkg_mux (sel : std_logic; one : ShiftCtrlEnum; zero : ShiftCtrlEnum) return ShiftCtrlEnum;
  subtype ShiftCtrlEnum_seq_type is std_logic_vector(1 downto 0);
  constant ShiftCtrlEnum_seq_DISABLE_1 : ShiftCtrlEnum_seq_type := "00";
  constant ShiftCtrlEnum_seq_SLL_1 : ShiftCtrlEnum_seq_type := "01";
  constant ShiftCtrlEnum_seq_SRL_1 : ShiftCtrlEnum_seq_type := "10";
  constant ShiftCtrlEnum_seq_SRA_1 : ShiftCtrlEnum_seq_type := "11";

  function pkg_mux (sel : std_logic; one : AluBitwiseCtrlEnum; zero : AluBitwiseCtrlEnum) return AluBitwiseCtrlEnum;
  subtype AluBitwiseCtrlEnum_seq_type is std_logic_vector(1 downto 0);
  constant AluBitwiseCtrlEnum_seq_XOR_1 : AluBitwiseCtrlEnum_seq_type := "00";
  constant AluBitwiseCtrlEnum_seq_OR_1 : AluBitwiseCtrlEnum_seq_type := "01";
  constant AluBitwiseCtrlEnum_seq_AND_1 : AluBitwiseCtrlEnum_seq_type := "10";

  function pkg_mux (sel : std_logic; one : Src2CtrlEnum; zero : Src2CtrlEnum) return Src2CtrlEnum;
  subtype Src2CtrlEnum_seq_type is std_logic_vector(1 downto 0);
  constant Src2CtrlEnum_seq_RS : Src2CtrlEnum_seq_type := "00";
  constant Src2CtrlEnum_seq_IMI : Src2CtrlEnum_seq_type := "01";
  constant Src2CtrlEnum_seq_IMS : Src2CtrlEnum_seq_type := "10";
  constant Src2CtrlEnum_seq_PC : Src2CtrlEnum_seq_type := "11";

  function pkg_mux (sel : std_logic; one : AluCtrlEnum; zero : AluCtrlEnum) return AluCtrlEnum;
  subtype AluCtrlEnum_seq_type is std_logic_vector(1 downto 0);
  constant AluCtrlEnum_seq_ADD_SUB : AluCtrlEnum_seq_type := "00";
  constant AluCtrlEnum_seq_SLT_SLTU : AluCtrlEnum_seq_type := "01";
  constant AluCtrlEnum_seq_BITWISE : AluCtrlEnum_seq_type := "10";

  function pkg_mux (sel : std_logic; one : Src1CtrlEnum; zero : Src1CtrlEnum) return Src1CtrlEnum;
  subtype Src1CtrlEnum_seq_type is std_logic_vector(1 downto 0);
  constant Src1CtrlEnum_seq_RS : Src1CtrlEnum_seq_type := "00";
  constant Src1CtrlEnum_seq_IMU : Src1CtrlEnum_seq_type := "01";
  constant Src1CtrlEnum_seq_PC_INCREMENT : Src1CtrlEnum_seq_type := "10";
  constant Src1CtrlEnum_seq_URS1 : Src1CtrlEnum_seq_type := "11";

end pkg_enum;

package body pkg_enum is
  function pkg_mux (sel : std_logic; one : Axi4ToApb3BridgePhase; zero : Axi4ToApb3BridgePhase) return Axi4ToApb3BridgePhase is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_toAxi4ToApb3BridgePhase_native (value : std_logic_vector(1 downto 0)) return Axi4ToApb3BridgePhase is
  begin
    case value is
      when "00" => return SETUP;
      when "01" => return ACCESS_1;
      when "10" => return RESPONSE;
      when others => return SETUP;
    end case;
  end;
  function pkg_toStdLogicVector_native (value : Axi4ToApb3BridgePhase) return std_logic_vector is
  begin
    case value is
      when SETUP => return "00";
      when ACCESS_1 => return "01";
      when RESPONSE => return "10";
      when others => return "00";
    end case;
  end;
  function pkg_mux (sel : std_logic; one : UartStopType; zero : UartStopType) return UartStopType is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : UartParityType; zero : UartParityType) return UartParityType is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : UartCtrlTxState; zero : UartCtrlTxState) return UartCtrlTxState is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_toUartCtrlTxState_native (value : std_logic_vector(2 downto 0)) return UartCtrlTxState is
  begin
    case value is
      when "000" => return IDLE;
      when "001" => return START;
      when "010" => return DATA;
      when "011" => return PARITY;
      when "100" => return STOP;
      when others => return IDLE;
    end case;
  end;
  function pkg_toStdLogicVector_native (value : UartCtrlTxState) return std_logic_vector is
  begin
    case value is
      when IDLE => return "000";
      when START => return "001";
      when DATA => return "010";
      when PARITY => return "011";
      when STOP => return "100";
      when others => return "000";
    end case;
  end;
  function pkg_mux (sel : std_logic; one : UartCtrlRxState; zero : UartCtrlRxState) return UartCtrlRxState is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_toUartCtrlRxState_native (value : std_logic_vector(2 downto 0)) return UartCtrlRxState is
  begin
    case value is
      when "000" => return IDLE;
      when "001" => return START;
      when "010" => return DATA;
      when "011" => return PARITY;
      when "100" => return STOP;
      when others => return IDLE;
    end case;
  end;
  function pkg_toStdLogicVector_native (value : UartCtrlRxState) return std_logic_vector is
  begin
    case value is
      when IDLE => return "000";
      when START => return "001";
      when DATA => return "010";
      when PARITY => return "011";
      when STOP => return "100";
      when others => return "000";
    end case;
  end;
  function pkg_mux (sel : std_logic; one : EnvCtrlEnum; zero : EnvCtrlEnum) return EnvCtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : BranchCtrlEnum; zero : BranchCtrlEnum) return BranchCtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : ShiftCtrlEnum; zero : ShiftCtrlEnum) return ShiftCtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : AluBitwiseCtrlEnum; zero : AluBitwiseCtrlEnum) return AluBitwiseCtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : Src2CtrlEnum; zero : Src2CtrlEnum) return Src2CtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : AluCtrlEnum; zero : AluCtrlEnum) return AluCtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : Src1CtrlEnum; zero : Src1CtrlEnum) return Src1CtrlEnum is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

end pkg_enum;


library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package pkg_scala2hdl is
  function pkg_extract (that : std_logic_vector; bitId : integer) return std_logic;
  function pkg_extract (that : std_logic_vector; base : unsigned; size : integer) return std_logic_vector;
  function pkg_cat (a : std_logic_vector; b : std_logic_vector) return std_logic_vector;
  function pkg_not (value : std_logic_vector) return std_logic_vector;
  function pkg_extract (that : unsigned; bitId : integer) return std_logic;
  function pkg_extract (that : unsigned; base : unsigned; size : integer) return unsigned;
  function pkg_cat (a : unsigned; b : unsigned) return unsigned;
  function pkg_not (value : unsigned) return unsigned;
  function pkg_extract (that : signed; bitId : integer) return std_logic;
  function pkg_extract (that : signed; base : unsigned; size : integer) return signed;
  function pkg_cat (a : signed; b : signed) return signed;
  function pkg_not (value : signed) return signed;

  function pkg_mux (sel : std_logic; one : std_logic; zero : std_logic) return std_logic;
  function pkg_mux (sel : std_logic; one : std_logic_vector; zero : std_logic_vector) return std_logic_vector;
  function pkg_mux (sel : std_logic; one : unsigned; zero : unsigned) return unsigned;
  function pkg_mux (sel : std_logic; one : signed; zero : signed) return signed;

  function pkg_toStdLogic (value : boolean) return std_logic;
  function pkg_toStdLogicVector (value : std_logic) return std_logic_vector;
  function pkg_toUnsigned (value : std_logic) return unsigned;
  function pkg_toSigned (value : std_logic) return signed;
  function pkg_stdLogicVector (lit : std_logic_vector) return std_logic_vector;
  function pkg_unsigned (lit : unsigned) return unsigned;
  function pkg_signed (lit : signed) return signed;

  function pkg_resize (that : std_logic_vector; width : integer) return std_logic_vector;
  function pkg_resize (that : unsigned; width : integer) return unsigned;
  function pkg_resize (that : signed; width : integer) return signed;

  function pkg_extract (that : std_logic_vector; high : integer; low : integer) return std_logic_vector;
  function pkg_extract (that : unsigned; high : integer; low : integer) return unsigned;
  function pkg_extract (that : signed; high : integer; low : integer) return signed;

  function pkg_shiftRight (that : std_logic_vector; size : natural) return std_logic_vector;
  function pkg_shiftRight (that : std_logic_vector; size : unsigned) return std_logic_vector;
  function pkg_shiftLeft (that : std_logic_vector; size : natural) return std_logic_vector;
  function pkg_shiftLeft (that : std_logic_vector; size : unsigned) return std_logic_vector;

  function pkg_shiftRight (that : unsigned; size : natural) return unsigned;
  function pkg_shiftRight (that : unsigned; size : unsigned) return unsigned;
  function pkg_shiftLeft (that : unsigned; size : natural) return unsigned;
  function pkg_shiftLeft (that : unsigned; size : unsigned) return unsigned;

  function pkg_shiftRight (that : signed; size : natural) return signed;
  function pkg_shiftRight (that : signed; size : unsigned) return signed;
  function pkg_shiftLeft (that : signed; size : natural) return signed;
  function pkg_shiftLeft (that : signed; size : unsigned; w : integer) return signed;

  function pkg_rotateLeft (that : std_logic_vector; size : unsigned) return std_logic_vector;
end  pkg_scala2hdl;

package body pkg_scala2hdl is
  function pkg_extract (that : std_logic_vector; bitId : integer) return std_logic is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : std_logic_vector; base : unsigned; size : integer) return std_logic_vector is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of std_logic_vector(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : std_logic_vector; b : std_logic_vector) return std_logic_vector is
    variable cat : std_logic_vector(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : std_logic_vector) return std_logic_vector is
    variable ret : std_logic_vector(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;

  function pkg_extract (that : unsigned; bitId : integer) return std_logic is
    alias temp : unsigned(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : unsigned; base : unsigned; size : integer) return unsigned is
    alias temp : unsigned(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of unsigned(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : unsigned; b : unsigned) return unsigned is
    variable cat : unsigned(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : unsigned) return unsigned is
    variable ret : unsigned(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;

  function pkg_extract (that : signed; bitId : integer) return std_logic is
    alias temp : signed(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : signed; base : unsigned; size : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of signed(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : signed; b : signed) return signed is
    variable cat : signed(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : signed) return signed is
    variable ret : signed(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;


  -- unsigned shifts
  function pkg_shiftRight (that : unsigned; size : natural) return unsigned is
    variable ret : unsigned(that'length-1 downto 0);
  begin
    if size >= that'length then
      return "";
    else
      ret := shift_right(that,size);
      return ret(that'length-1-size downto 0);
    end if;
  end pkg_shiftRight;

  function pkg_shiftRight (that : unsigned; size : unsigned) return unsigned is
    variable ret : unsigned(that'length-1 downto 0);
  begin
    ret := shift_right(that,to_integer(size));
    return ret;
  end pkg_shiftRight;

  function pkg_shiftLeft (that : unsigned; size : natural) return unsigned is
  begin
    return shift_left(resize(that,that'length + size),size);
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : unsigned; size : unsigned) return unsigned is
  begin
    return shift_left(resize(that,that'length + 2**size'length - 1),to_integer(size));
  end pkg_shiftLeft;

  -- std_logic_vector shifts
  function pkg_shiftRight (that : std_logic_vector; size : natural) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftRight (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftLeft (that : std_logic_vector; size : natural) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  -- signed shifts
  function pkg_shiftRight (that : signed; size : natural) return signed is
  begin
    return signed(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftRight (that : signed; size : unsigned) return signed is
  begin
    return shift_right(that,to_integer(size));
  end pkg_shiftRight;

  function pkg_shiftLeft (that : signed; size : natural) return signed is
  begin
    return signed(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : signed; size : unsigned; w : integer) return signed is
  begin
    return shift_left(resize(that,w),to_integer(size));
  end pkg_shiftLeft;

  function pkg_rotateLeft (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(rotate_left(unsigned(that),to_integer(size)));
  end pkg_rotateLeft;

  function pkg_extract (that : std_logic_vector; high : integer; low : integer) return std_logic_vector is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_extract (that : unsigned; high : integer; low : integer) return unsigned is
    alias temp : unsigned(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_extract (that : signed; high : integer; low : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_mux (sel : std_logic; one : std_logic; zero : std_logic) return std_logic is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : std_logic_vector; zero : std_logic_vector) return std_logic_vector is
    variable ret : std_logic_vector(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : unsigned; zero : unsigned) return unsigned is
    variable ret : unsigned(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : signed; zero : signed) return signed is
    variable ret : signed(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_toStdLogic (value : boolean) return std_logic is
  begin
    if value = true then
      return '1';
    else
      return '0';
    end if;
  end pkg_toStdLogic;

  function pkg_toStdLogicVector (value : std_logic) return std_logic_vector is
    variable ret : std_logic_vector(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toStdLogicVector;

  function pkg_toUnsigned (value : std_logic) return unsigned is
    variable ret : unsigned(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toUnsigned;

  function pkg_toSigned (value : std_logic) return signed is
    variable ret : signed(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toSigned;

  function pkg_stdLogicVector (lit : std_logic_vector) return std_logic_vector is
    alias ret : std_logic_vector(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_stdLogicVector;

  function pkg_unsigned (lit : unsigned) return unsigned is
    alias ret : unsigned(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_unsigned;

  function pkg_signed (lit : signed) return signed is
    alias ret : signed(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_signed;

  function pkg_resize (that : std_logic_vector; width : integer) return std_logic_vector is
  begin
    return std_logic_vector(resize(unsigned(that),width));
  end pkg_resize;

  function pkg_resize (that : unsigned; width : integer) return unsigned is
    variable ret : unsigned(width-1 downto 0);
  begin
    if that'length = 0 then
       ret := (others => '0');
    else
       ret := resize(that,width);
    end if;
    return ret;
  end pkg_resize;
  function pkg_resize (that : signed; width : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;
    variable ret : signed(width-1 downto 0);
  begin
    if temp'length = 0 then
       ret := (others => '0');
    elsif temp'length >= width then
       ret := temp(width-1 downto 0);
    else
       ret := resize(temp,width);
    end if;
    return ret;
  end pkg_resize;
end pkg_scala2hdl;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity BufferCC is
  port(
    io_dataIn : in std_logic;
    io_dataOut : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end BufferCC;

architecture arch of BufferCC is
  attribute async_reg : string;

  signal buffers_0 : std_logic;
  attribute async_reg of buffers_0 : signal is "true";
  signal buffers_1 : std_logic;
  attribute async_reg of buffers_1 : signal is "true";
begin
  io_dataOut <= buffers_1;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      buffers_0 <= pkg_toStdLogic(false);
      buffers_1 <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity UartCtrlTx is
  port(
    io_configFrame_dataLength : in unsigned(2 downto 0);
    io_configFrame_stop : in UartStopType_seq_type;
    io_configFrame_parity : in UartParityType_seq_type;
    io_samplingTick : in std_logic;
    io_write_valid : in std_logic;
    io_write_ready : out std_logic;
    io_write_payload : in std_logic_vector(7 downto 0);
    io_cts : in std_logic;
    io_txd : out std_logic;
    io_break : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end UartCtrlTx;

architecture arch of UartCtrlTx is

  signal clockDivider_counter_willIncrement : std_logic;
  signal clockDivider_counter_willClear : std_logic;
  signal clockDivider_counter_valueNext : unsigned(2 downto 0);
  signal clockDivider_counter_value : unsigned(2 downto 0);
  signal clockDivider_counter_willOverflowIfInc : std_logic;
  signal clockDivider_counter_willOverflow : std_logic;
  signal tickCounter_value : unsigned(2 downto 0);
  signal stateMachine_state : UartCtrlTxState;
  signal stateMachine_parity : std_logic;
  signal stateMachine_txd : std_logic;
  signal when_UartCtrlTx_l58 : std_logic;
  signal when_UartCtrlTx_l73 : std_logic;
  signal when_UartCtrlTx_l76 : std_logic;
  signal when_UartCtrlTx_l93 : std_logic;
  signal zz_io_txd : std_logic;
begin
  process(io_samplingTick)
  begin
    clockDivider_counter_willIncrement <= pkg_toStdLogic(false);
    if io_samplingTick = '1' then
      clockDivider_counter_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  clockDivider_counter_willClear <= pkg_toStdLogic(false);
  clockDivider_counter_willOverflowIfInc <= pkg_toStdLogic(clockDivider_counter_value = pkg_unsigned("100"));
  clockDivider_counter_willOverflow <= (clockDivider_counter_willOverflowIfInc and clockDivider_counter_willIncrement);
  process(clockDivider_counter_willOverflow,clockDivider_counter_value,clockDivider_counter_willIncrement,clockDivider_counter_willClear)
  begin
    if clockDivider_counter_willOverflow = '1' then
      clockDivider_counter_valueNext <= pkg_unsigned("000");
    else
      clockDivider_counter_valueNext <= (clockDivider_counter_value + pkg_resize(unsigned(pkg_toStdLogicVector(clockDivider_counter_willIncrement)),3));
    end if;
    if clockDivider_counter_willClear = '1' then
      clockDivider_counter_valueNext <= pkg_unsigned("000");
    end if;
  end process;

  process(stateMachine_state,io_write_payload,tickCounter_value,stateMachine_parity)
  begin
    stateMachine_txd <= pkg_toStdLogic(true);
    case stateMachine_state is
      when pkg_enum.IDLE =>
      when pkg_enum.START =>
        stateMachine_txd <= pkg_toStdLogic(false);
      when pkg_enum.DATA =>
        stateMachine_txd <= pkg_extract(io_write_payload,to_integer(tickCounter_value));
      when pkg_enum.PARITY =>
        stateMachine_txd <= stateMachine_parity;
      when others =>
    end case;
  end process;

  process(io_break,stateMachine_state,clockDivider_counter_willOverflow,when_UartCtrlTx_l73)
  begin
    io_write_ready <= io_break;
    case stateMachine_state is
      when pkg_enum.IDLE =>
      when pkg_enum.START =>
      when pkg_enum.DATA =>
        if clockDivider_counter_willOverflow = '1' then
          if when_UartCtrlTx_l73 = '1' then
            io_write_ready <= pkg_toStdLogic(true);
          end if;
        end if;
      when pkg_enum.PARITY =>
      when others =>
    end case;
  end process;

  when_UartCtrlTx_l58 <= ((io_write_valid and (not io_cts)) and clockDivider_counter_willOverflow);
  when_UartCtrlTx_l73 <= pkg_toStdLogic(tickCounter_value = io_configFrame_dataLength);
  when_UartCtrlTx_l76 <= pkg_toStdLogic(io_configFrame_parity = UartParityType_seq_NONE);
  when_UartCtrlTx_l93 <= pkg_toStdLogic(tickCounter_value = pkg_resize(pkg_mux(pkg_toStdLogic(io_configFrame_stop = UartStopType_seq_ONE),pkg_unsigned("0"),pkg_unsigned("1")),3));
  io_txd <= zz_io_txd;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      clockDivider_counter_value <= pkg_unsigned("000");
      stateMachine_state <= pkg_enum.IDLE;
      zz_io_txd <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      clockDivider_counter_value <= clockDivider_counter_valueNext;
      case stateMachine_state is
        when pkg_enum.IDLE =>
          if when_UartCtrlTx_l58 = '1' then
            stateMachine_state <= pkg_enum.START;
          end if;
        when pkg_enum.START =>
          if clockDivider_counter_willOverflow = '1' then
            stateMachine_state <= pkg_enum.DATA;
          end if;
        when pkg_enum.DATA =>
          if clockDivider_counter_willOverflow = '1' then
            if when_UartCtrlTx_l73 = '1' then
              if when_UartCtrlTx_l76 = '1' then
                stateMachine_state <= pkg_enum.STOP;
              else
                stateMachine_state <= pkg_enum.PARITY;
              end if;
            end if;
          end if;
        when pkg_enum.PARITY =>
          if clockDivider_counter_willOverflow = '1' then
            stateMachine_state <= pkg_enum.STOP;
          end if;
        when others =>
          if clockDivider_counter_willOverflow = '1' then
            if when_UartCtrlTx_l93 = '1' then
              stateMachine_state <= pkg_mux(io_write_valid,pkg_enum.START,pkg_enum.IDLE);
            end if;
          end if;
      end case;
      zz_io_txd <= (stateMachine_txd and (not io_break));
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if clockDivider_counter_willOverflow = '1' then
        tickCounter_value <= (tickCounter_value + pkg_unsigned("001"));
      end if;
      if clockDivider_counter_willOverflow = '1' then
        stateMachine_parity <= (stateMachine_parity xor stateMachine_txd);
      end if;
      case stateMachine_state is
        when pkg_enum.IDLE =>
        when pkg_enum.START =>
          if clockDivider_counter_willOverflow = '1' then
            stateMachine_parity <= pkg_toStdLogic(io_configFrame_parity = UartParityType_seq_ODD);
            tickCounter_value <= pkg_unsigned("000");
          end if;
        when pkg_enum.DATA =>
          if clockDivider_counter_willOverflow = '1' then
            if when_UartCtrlTx_l73 = '1' then
              tickCounter_value <= pkg_unsigned("000");
            end if;
          end if;
        when pkg_enum.PARITY =>
          if clockDivider_counter_willOverflow = '1' then
            tickCounter_value <= pkg_unsigned("000");
          end if;
        when others =>
      end case;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity UartCtrlRx is
  port(
    io_configFrame_dataLength : in unsigned(2 downto 0);
    io_configFrame_stop : in UartStopType_seq_type;
    io_configFrame_parity : in UartParityType_seq_type;
    io_samplingTick : in std_logic;
    io_read_valid : out std_logic;
    io_read_ready : in std_logic;
    io_read_payload : out std_logic_vector(7 downto 0);
    io_rxd : in std_logic;
    io_rts : out std_logic;
    io_error : out std_logic;
    io_break : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end UartCtrlRx;

architecture arch of UartCtrlRx is
  signal io_rxd_buffercc_io_dataOut : std_logic;

  signal zz_io_rts : std_logic;
  signal sampler_synchroniser : std_logic;
  signal sampler_samples_0 : std_logic;
  signal sampler_samples_1 : std_logic;
  signal sampler_samples_2 : std_logic;
  signal sampler_value : std_logic;
  signal sampler_tick : std_logic;
  signal bitTimer_counter : unsigned(2 downto 0);
  signal bitTimer_tick : std_logic;
  signal when_UartCtrlRx_l43 : std_logic;
  signal bitCounter_value : unsigned(2 downto 0);
  signal break_counter : unsigned(6 downto 0);
  signal break_valid : std_logic;
  signal when_UartCtrlRx_l69 : std_logic;
  signal stateMachine_state : UartCtrlRxState;
  signal stateMachine_parity : std_logic;
  signal stateMachine_shifter : std_logic_vector(7 downto 0);
  signal stateMachine_validReg : std_logic;
  signal when_UartCtrlRx_l93 : std_logic;
  signal when_UartCtrlRx_l103 : std_logic;
  signal when_UartCtrlRx_l111 : std_logic;
  signal when_UartCtrlRx_l113 : std_logic;
  signal when_UartCtrlRx_l125 : std_logic;
  signal when_UartCtrlRx_l136 : std_logic;
  signal when_UartCtrlRx_l139 : std_logic;
begin
  io_rxd_buffercc : entity work.BufferCC
    port map ( 
      io_dataIn => io_rxd,
      io_dataOut => io_rxd_buffercc_io_dataOut,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  process(stateMachine_state,bitTimer_tick,when_UartCtrlRx_l125,when_UartCtrlRx_l136)
  begin
    io_error <= pkg_toStdLogic(false);
    case stateMachine_state is
      when pkg_enum.IDLE =>
      when pkg_enum.START =>
      when pkg_enum.DATA =>
      when pkg_enum.PARITY =>
        if bitTimer_tick = '1' then
          if when_UartCtrlRx_l125 = '0' then
            io_error <= pkg_toStdLogic(true);
          end if;
        end if;
      when others =>
        if bitTimer_tick = '1' then
          if when_UartCtrlRx_l136 = '1' then
            io_error <= pkg_toStdLogic(true);
          end if;
        end if;
    end case;
  end process;

  io_rts <= zz_io_rts;
  sampler_synchroniser <= io_rxd_buffercc_io_dataOut;
  sampler_samples_0 <= sampler_synchroniser;
  process(sampler_tick,when_UartCtrlRx_l43)
  begin
    bitTimer_tick <= pkg_toStdLogic(false);
    if sampler_tick = '1' then
      if when_UartCtrlRx_l43 = '1' then
        bitTimer_tick <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  when_UartCtrlRx_l43 <= pkg_toStdLogic(bitTimer_counter = pkg_unsigned("000"));
  break_valid <= pkg_toStdLogic(break_counter = pkg_unsigned("1000001"));
  when_UartCtrlRx_l69 <= (io_samplingTick and (not break_valid));
  io_break <= break_valid;
  io_read_valid <= stateMachine_validReg;
  when_UartCtrlRx_l93 <= ((sampler_tick and (not sampler_value)) and (not break_valid));
  when_UartCtrlRx_l103 <= pkg_toStdLogic(sampler_value = pkg_toStdLogic(true));
  when_UartCtrlRx_l111 <= pkg_toStdLogic(bitCounter_value = io_configFrame_dataLength);
  when_UartCtrlRx_l113 <= pkg_toStdLogic(io_configFrame_parity = UartParityType_seq_NONE);
  when_UartCtrlRx_l125 <= pkg_toStdLogic(stateMachine_parity = sampler_value);
  when_UartCtrlRx_l136 <= (not sampler_value);
  when_UartCtrlRx_l139 <= pkg_toStdLogic(bitCounter_value = pkg_resize(pkg_mux(pkg_toStdLogic(io_configFrame_stop = UartStopType_seq_ONE),pkg_unsigned("0"),pkg_unsigned("1")),3));
  io_read_payload <= stateMachine_shifter;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      zz_io_rts <= pkg_toStdLogic(false);
      sampler_samples_1 <= pkg_toStdLogic(true);
      sampler_samples_2 <= pkg_toStdLogic(true);
      sampler_value <= pkg_toStdLogic(true);
      sampler_tick <= pkg_toStdLogic(false);
      break_counter <= pkg_unsigned("0000000");
      stateMachine_state <= pkg_enum.IDLE;
      stateMachine_validReg <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      zz_io_rts <= (not io_read_ready);
      if io_samplingTick = '1' then
        sampler_samples_1 <= sampler_samples_0;
      end if;
      if io_samplingTick = '1' then
        sampler_samples_2 <= sampler_samples_1;
      end if;
      sampler_value <= (((pkg_toStdLogic(false) or ((pkg_toStdLogic(true) and sampler_samples_0) and sampler_samples_1)) or ((pkg_toStdLogic(true) and sampler_samples_0) and sampler_samples_2)) or ((pkg_toStdLogic(true) and sampler_samples_1) and sampler_samples_2));
      sampler_tick <= io_samplingTick;
      if sampler_value = '1' then
        break_counter <= pkg_unsigned("0000000");
      else
        if when_UartCtrlRx_l69 = '1' then
          break_counter <= (break_counter + pkg_unsigned("0000001"));
        end if;
      end if;
      stateMachine_validReg <= pkg_toStdLogic(false);
      case stateMachine_state is
        when pkg_enum.IDLE =>
          if when_UartCtrlRx_l93 = '1' then
            stateMachine_state <= pkg_enum.START;
          end if;
        when pkg_enum.START =>
          if bitTimer_tick = '1' then
            stateMachine_state <= pkg_enum.DATA;
            if when_UartCtrlRx_l103 = '1' then
              stateMachine_state <= pkg_enum.IDLE;
            end if;
          end if;
        when pkg_enum.DATA =>
          if bitTimer_tick = '1' then
            if when_UartCtrlRx_l111 = '1' then
              if when_UartCtrlRx_l113 = '1' then
                stateMachine_state <= pkg_enum.STOP;
                stateMachine_validReg <= pkg_toStdLogic(true);
              else
                stateMachine_state <= pkg_enum.PARITY;
              end if;
            end if;
          end if;
        when pkg_enum.PARITY =>
          if bitTimer_tick = '1' then
            if when_UartCtrlRx_l125 = '1' then
              stateMachine_state <= pkg_enum.STOP;
              stateMachine_validReg <= pkg_toStdLogic(true);
            else
              stateMachine_state <= pkg_enum.IDLE;
            end if;
          end if;
        when others =>
          if bitTimer_tick = '1' then
            if when_UartCtrlRx_l136 = '1' then
              stateMachine_state <= pkg_enum.IDLE;
            else
              if when_UartCtrlRx_l139 = '1' then
                stateMachine_state <= pkg_enum.IDLE;
              end if;
            end if;
          end if;
      end case;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if sampler_tick = '1' then
        bitTimer_counter <= (bitTimer_counter - pkg_unsigned("001"));
        if when_UartCtrlRx_l43 = '1' then
          bitTimer_counter <= pkg_unsigned("100");
        end if;
      end if;
      if bitTimer_tick = '1' then
        bitCounter_value <= (bitCounter_value + pkg_unsigned("001"));
      end if;
      if bitTimer_tick = '1' then
        stateMachine_parity <= (stateMachine_parity xor sampler_value);
      end if;
      case stateMachine_state is
        when pkg_enum.IDLE =>
          if when_UartCtrlRx_l93 = '1' then
            bitTimer_counter <= pkg_unsigned("001");
          end if;
        when pkg_enum.START =>
          if bitTimer_tick = '1' then
            bitCounter_value <= pkg_unsigned("000");
            stateMachine_parity <= pkg_toStdLogic(io_configFrame_parity = UartParityType_seq_ODD);
          end if;
        when pkg_enum.DATA =>
          if bitTimer_tick = '1' then
            stateMachine_shifter(to_integer(bitCounter_value)) <= sampler_value;
            if when_UartCtrlRx_l111 = '1' then
              bitCounter_value <= pkg_unsigned("000");
            end if;
          end if;
        when pkg_enum.PARITY =>
          if bitTimer_tick = '1' then
            bitCounter_value <= pkg_unsigned("000");
          end if;
        when others =>
      end case;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity BufferCC_1 is
  port(
    io_dataIn : in std_logic;
    io_dataOut : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_systemReset : in std_logic
  );
end BufferCC_1;

architecture arch of BufferCC_1 is
  attribute async_reg : string;

  signal buffers_0 : std_logic;
  attribute async_reg of buffers_0 : signal is "true";
  signal buffers_1 : std_logic;
  attribute async_reg of buffers_1 : signal is "true";
begin
  io_dataOut <= buffers_1;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity BufferCC_2 is
  port(
    io_dataIn : in std_logic_vector(31 downto 0);
    io_dataOut : out std_logic_vector(31 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end BufferCC_2;

architecture arch of BufferCC_2 is
  attribute async_reg : string;

  signal buffers_0 : std_logic_vector(31 downto 0);
  attribute async_reg of buffers_0 : signal is "true";
  signal buffers_1 : std_logic_vector(31 downto 0);
  attribute async_reg of buffers_1 : signal is "true";
begin
  io_dataOut <= buffers_1;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity UartCtrl is
  port(
    io_config_frame_dataLength : in unsigned(2 downto 0);
    io_config_frame_stop : in UartStopType_seq_type;
    io_config_frame_parity : in UartParityType_seq_type;
    io_config_clockDivider : in unsigned(19 downto 0);
    io_write_valid : in std_logic;
    io_write_ready : out std_logic;
    io_write_payload : in std_logic_vector(7 downto 0);
    io_read_valid : out std_logic;
    io_read_ready : in std_logic;
    io_read_payload : out std_logic_vector(7 downto 0);
    io_uart_txd : out std_logic;
    io_uart_rxd : in std_logic;
    io_readError : out std_logic;
    io_writeBreak : in std_logic;
    io_readBreak : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end UartCtrl;

architecture arch of UartCtrl is
  signal tx_io_write_ready : std_logic;
  signal tx_io_txd : std_logic;
  signal rx_io_read_valid : std_logic;
  signal rx_io_read_payload : std_logic_vector(7 downto 0);
  signal rx_io_rts : std_logic;
  signal rx_io_error : std_logic;
  signal rx_io_break : std_logic;

  signal clockDivider_counter : unsigned(19 downto 0);
  signal clockDivider_tick : std_logic;
  signal clockDivider_tickReg : std_logic;
  signal io_write_thrown_valid : std_logic;
  signal io_write_thrown_ready : std_logic;
  signal io_write_thrown_payload : std_logic_vector(7 downto 0);
begin
  tx : entity work.UartCtrlTx
    port map ( 
      io_configFrame_dataLength => io_config_frame_dataLength,
      io_configFrame_stop => io_config_frame_stop,
      io_configFrame_parity => io_config_frame_parity,
      io_samplingTick => clockDivider_tickReg,
      io_write_valid => io_write_thrown_valid,
      io_write_ready => tx_io_write_ready,
      io_write_payload => io_write_thrown_payload,
      io_cts => pkg_toStdLogic(false),
      io_txd => tx_io_txd,
      io_break => io_writeBreak,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  rx : entity work.UartCtrlRx
    port map ( 
      io_configFrame_dataLength => io_config_frame_dataLength,
      io_configFrame_stop => io_config_frame_stop,
      io_configFrame_parity => io_config_frame_parity,
      io_samplingTick => clockDivider_tickReg,
      io_read_valid => rx_io_read_valid,
      io_read_ready => io_read_ready,
      io_read_payload => rx_io_read_payload,
      io_rxd => io_uart_rxd,
      io_rts => rx_io_rts,
      io_error => rx_io_error,
      io_break => rx_io_break,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  clockDivider_tick <= pkg_toStdLogic(clockDivider_counter = pkg_unsigned("00000000000000000000"));
  process(io_write_valid,rx_io_break)
  begin
    io_write_thrown_valid <= io_write_valid;
    if rx_io_break = '1' then
      io_write_thrown_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  process(io_write_thrown_ready,rx_io_break)
  begin
    io_write_ready <= io_write_thrown_ready;
    if rx_io_break = '1' then
      io_write_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  io_write_thrown_payload <= io_write_payload;
  io_write_thrown_ready <= tx_io_write_ready;
  io_read_valid <= rx_io_read_valid;
  io_read_payload <= rx_io_read_payload;
  io_uart_txd <= tx_io_txd;
  io_readError <= rx_io_error;
  io_readBreak <= rx_io_break;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      clockDivider_counter <= pkg_unsigned("00000000000000000000");
      clockDivider_tickReg <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      clockDivider_tickReg <= clockDivider_tick;
      clockDivider_counter <= (clockDivider_counter - pkg_unsigned("00000000000000000001"));
      if clockDivider_tick = '1' then
        clockDivider_counter <= io_config_clockDivider;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamFifo is
  port(
    io_push_valid : in std_logic;
    io_push_ready : out std_logic;
    io_push_payload : in std_logic_vector(7 downto 0);
    io_pop_valid : out std_logic;
    io_pop_ready : in std_logic;
    io_pop_payload : out std_logic_vector(7 downto 0);
    io_flush : in std_logic;
    io_occupancy : out unsigned(4 downto 0);
    io_availability : out unsigned(4 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamFifo;

architecture arch of StreamFifo is
  signal zz_logic_ram_port0 : std_logic_vector(7 downto 0);
  signal io_push_ready_read_buffer : std_logic;
  signal io_pop_valid_read_buffer : std_logic;
  signal zz_logic_ram_port : std_logic;
  signal zz_io_pop_payload : std_logic;

  signal zz_1 : std_logic;
  signal logic_pushPtr_willIncrement : std_logic;
  signal logic_pushPtr_willClear : std_logic;
  signal logic_pushPtr_valueNext : unsigned(3 downto 0);
  signal logic_pushPtr_value : unsigned(3 downto 0);
  signal logic_pushPtr_willOverflowIfInc : std_logic;
  signal logic_pushPtr_willOverflow : std_logic;
  signal logic_popPtr_willIncrement : std_logic;
  signal logic_popPtr_willClear : std_logic;
  signal logic_popPtr_valueNext : unsigned(3 downto 0);
  signal logic_popPtr_value : unsigned(3 downto 0);
  signal logic_popPtr_willOverflowIfInc : std_logic;
  signal logic_popPtr_willOverflow : std_logic;
  signal logic_ptrMatch : std_logic;
  signal logic_risingOccupancy : std_logic;
  signal logic_pushing : std_logic;
  signal logic_popping : std_logic;
  signal logic_empty : std_logic;
  signal logic_full : std_logic;
  signal zz_io_pop_valid : std_logic;
  signal when_Stream_l946 : std_logic;
  signal logic_ptrDif : unsigned(3 downto 0);
  type logic_ram_type is array (0 to 15) of std_logic_vector(7 downto 0);
  signal logic_ram : logic_ram_type;
begin
  io_push_ready <= io_push_ready_read_buffer;
  io_pop_valid <= io_pop_valid_read_buffer;
  zz_io_pop_payload <= pkg_toStdLogic(true);
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_io_pop_payload = '1' then
        zz_logic_ram_port0 <= logic_ram(to_integer(logic_popPtr_valueNext));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_1 = '1' then
        logic_ram(to_integer(logic_pushPtr_value)) <= io_push_payload;
      end if;
    end if;
  end process;

  process(logic_pushing)
  begin
    zz_1 <= pkg_toStdLogic(false);
    if logic_pushing = '1' then
      zz_1 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(logic_pushing)
  begin
    logic_pushPtr_willIncrement <= pkg_toStdLogic(false);
    if logic_pushing = '1' then
      logic_pushPtr_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_flush)
  begin
    logic_pushPtr_willClear <= pkg_toStdLogic(false);
    if io_flush = '1' then
      logic_pushPtr_willClear <= pkg_toStdLogic(true);
    end if;
  end process;

  logic_pushPtr_willOverflowIfInc <= pkg_toStdLogic(logic_pushPtr_value = pkg_unsigned("1111"));
  logic_pushPtr_willOverflow <= (logic_pushPtr_willOverflowIfInc and logic_pushPtr_willIncrement);
  process(logic_pushPtr_value,logic_pushPtr_willIncrement,logic_pushPtr_willClear)
  begin
    logic_pushPtr_valueNext <= (logic_pushPtr_value + pkg_resize(unsigned(pkg_toStdLogicVector(logic_pushPtr_willIncrement)),4));
    if logic_pushPtr_willClear = '1' then
      logic_pushPtr_valueNext <= pkg_unsigned("0000");
    end if;
  end process;

  process(logic_popping)
  begin
    logic_popPtr_willIncrement <= pkg_toStdLogic(false);
    if logic_popping = '1' then
      logic_popPtr_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_flush)
  begin
    logic_popPtr_willClear <= pkg_toStdLogic(false);
    if io_flush = '1' then
      logic_popPtr_willClear <= pkg_toStdLogic(true);
    end if;
  end process;

  logic_popPtr_willOverflowIfInc <= pkg_toStdLogic(logic_popPtr_value = pkg_unsigned("1111"));
  logic_popPtr_willOverflow <= (logic_popPtr_willOverflowIfInc and logic_popPtr_willIncrement);
  process(logic_popPtr_value,logic_popPtr_willIncrement,logic_popPtr_willClear)
  begin
    logic_popPtr_valueNext <= (logic_popPtr_value + pkg_resize(unsigned(pkg_toStdLogicVector(logic_popPtr_willIncrement)),4));
    if logic_popPtr_willClear = '1' then
      logic_popPtr_valueNext <= pkg_unsigned("0000");
    end if;
  end process;

  logic_ptrMatch <= pkg_toStdLogic(logic_pushPtr_value = logic_popPtr_value);
  logic_pushing <= (io_push_valid and io_push_ready_read_buffer);
  logic_popping <= (io_pop_valid_read_buffer and io_pop_ready);
  logic_empty <= (logic_ptrMatch and (not logic_risingOccupancy));
  logic_full <= (logic_ptrMatch and logic_risingOccupancy);
  io_push_ready_read_buffer <= (not logic_full);
  io_pop_valid_read_buffer <= ((not logic_empty) and (not (zz_io_pop_valid and (not logic_full))));
  io_pop_payload <= zz_logic_ram_port0;
  when_Stream_l946 <= pkg_toStdLogic(logic_pushing /= logic_popping);
  logic_ptrDif <= (logic_pushPtr_value - logic_popPtr_value);
  io_occupancy <= unsigned(pkg_cat(pkg_toStdLogicVector((logic_risingOccupancy and logic_ptrMatch)),std_logic_vector(logic_ptrDif)));
  io_availability <= unsigned(pkg_cat(pkg_toStdLogicVector(((not logic_risingOccupancy) and logic_ptrMatch)),std_logic_vector((logic_popPtr_value - logic_pushPtr_value))));
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      logic_pushPtr_value <= pkg_unsigned("0000");
      logic_popPtr_value <= pkg_unsigned("0000");
      logic_risingOccupancy <= pkg_toStdLogic(false);
      zz_io_pop_valid <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      zz_io_pop_valid <= pkg_toStdLogic(logic_popPtr_valueNext = logic_pushPtr_value);
      if when_Stream_l946 = '1' then
        logic_risingOccupancy <= logic_pushing;
      end if;
      if io_flush = '1' then
        logic_risingOccupancy <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

end arch;


--StreamFifo_1 replaced by StreamFifo

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Prescaler is
  port(
    io_clear : in std_logic;
    io_limit : in unsigned(31 downto 0);
    io_overflow : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Prescaler;

architecture arch of Prescaler is
  signal io_overflow_read_buffer : std_logic;

  signal counter : unsigned(31 downto 0);
  signal when_Prescaler_l17 : std_logic;
begin
  io_overflow <= io_overflow_read_buffer;
  when_Prescaler_l17 <= (io_clear or io_overflow_read_buffer);
  io_overflow_read_buffer <= pkg_toStdLogic(counter = io_limit);
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      counter <= (counter + pkg_unsigned("00000000000000000000000000000001"));
      if when_Prescaler_l17 = '1' then
        counter <= pkg_unsigned("00000000000000000000000000000000");
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Timer is
  port(
    io_tick : in std_logic;
    io_clear : in std_logic;
    io_limit : in unsigned(15 downto 0);
    io_full : out std_logic;
    io_value : out unsigned(15 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Timer;

architecture arch of Timer is

  signal counter : unsigned(15 downto 0);
  signal limitHit : std_logic;
  signal inhibitFull : std_logic;
begin
  limitHit <= pkg_toStdLogic(counter = io_limit);
  io_full <= ((limitHit and io_tick) and (not inhibitFull));
  io_value <= counter;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      inhibitFull <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if io_tick = '1' then
        inhibitFull <= limitHit;
      end if;
      if io_clear = '1' then
        inhibitFull <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_tick = '1' then
        counter <= (counter + pkg_resize(unsigned(pkg_toStdLogicVector((not limitHit))),16));
      end if;
      if io_clear = '1' then
        counter <= pkg_unsigned("0000000000000000");
      end if;
    end if;
  end process;

end arch;


--Timer_1 replaced by Timer

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity InterruptCtrl is
  port(
    io_inputs : in std_logic_vector(1 downto 0);
    io_clears : in std_logic_vector(1 downto 0);
    io_masks : in std_logic_vector(1 downto 0);
    io_pendings : out std_logic_vector(1 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end InterruptCtrl;

architecture arch of InterruptCtrl is

  signal pendings : std_logic_vector(1 downto 0);
begin
  io_pendings <= (pendings and io_masks);
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      pendings <= pkg_stdLogicVector("00");
    elsif rising_edge(io_mainClk) then
      pendings <= ((pendings and pkg_not(io_clears)) or io_inputs);
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity InstructionCache is
  port(
    io_flush : in std_logic;
    io_cpu_prefetch_isValid : in std_logic;
    io_cpu_prefetch_haltIt : out std_logic;
    io_cpu_prefetch_pc : in unsigned(31 downto 0);
    io_cpu_fetch_isValid : in std_logic;
    io_cpu_fetch_isStuck : in std_logic;
    io_cpu_fetch_isRemoved : in std_logic;
    io_cpu_fetch_pc : in unsigned(31 downto 0);
    io_cpu_fetch_data : out std_logic_vector(31 downto 0);
    io_cpu_fetch_mmuRsp_physicalAddress : in unsigned(31 downto 0);
    io_cpu_fetch_mmuRsp_isIoAccess : in std_logic;
    io_cpu_fetch_mmuRsp_isPaging : in std_logic;
    io_cpu_fetch_mmuRsp_allowRead : in std_logic;
    io_cpu_fetch_mmuRsp_allowWrite : in std_logic;
    io_cpu_fetch_mmuRsp_allowExecute : in std_logic;
    io_cpu_fetch_mmuRsp_exception : in std_logic;
    io_cpu_fetch_mmuRsp_refilling : in std_logic;
    io_cpu_fetch_mmuRsp_bypassTranslation : in std_logic;
    io_cpu_fetch_physicalAddress : out unsigned(31 downto 0);
    io_cpu_decode_isValid : in std_logic;
    io_cpu_decode_isStuck : in std_logic;
    io_cpu_decode_pc : in unsigned(31 downto 0);
    io_cpu_decode_physicalAddress : out unsigned(31 downto 0);
    io_cpu_decode_data : out std_logic_vector(31 downto 0);
    io_cpu_decode_cacheMiss : out std_logic;
    io_cpu_decode_error : out std_logic;
    io_cpu_decode_mmuRefilling : out std_logic;
    io_cpu_decode_mmuException : out std_logic;
    io_cpu_decode_isUser : in std_logic;
    io_cpu_fill_valid : in std_logic;
    io_cpu_fill_payload : in unsigned(31 downto 0);
    io_mem_cmd_valid : out std_logic;
    io_mem_cmd_ready : in std_logic;
    io_mem_cmd_payload_address : out unsigned(31 downto 0);
    io_mem_cmd_payload_size : out unsigned(2 downto 0);
    io_mem_rsp_valid : in std_logic;
    io_mem_rsp_payload_data : in std_logic_vector(31 downto 0);
    io_mem_rsp_payload_error : in std_logic;
    zz_when_Fetcher_l398 : in unsigned(2 downto 0);
    zz_io_cpu_fetch_data_regNextWhen : in std_logic_vector(31 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end InstructionCache;

architecture arch of InstructionCache is
  signal zz_banks_0_port0 : std_logic_vector(31 downto 0);
  signal zz_ways_0_tags_port0 : std_logic_vector(20 downto 0);
  signal io_mem_cmd_valid_read_buffer : std_logic;
  signal io_cpu_fetch_data_read_buffer : std_logic_vector(31 downto 0);
  signal zz_ways_0_tags_port : std_logic_vector(20 downto 0);
  attribute keep : boolean;
  attribute syn_keep : boolean;

  signal zz_1 : std_logic;
  signal zz_2 : std_logic;
  signal lineLoader_fire : std_logic;
  signal lineLoader_valid : std_logic;
  signal lineLoader_address : unsigned(31 downto 0);
  attribute keep of lineLoader_address : signal is true;
  attribute syn_keep of lineLoader_address : signal is true;
  signal lineLoader_hadError : std_logic;
  signal lineLoader_flushPending : std_logic;
  signal lineLoader_flushCounter : unsigned(8 downto 0);
  signal when_InstructionCache_l338 : std_logic;
  signal zz_when_InstructionCache_l342 : std_logic;
  signal when_InstructionCache_l342 : std_logic;
  signal when_InstructionCache_l351 : std_logic;
  signal lineLoader_cmdSent : std_logic;
  signal io_mem_cmd_fire : std_logic;
  signal when_Utils_l485 : std_logic;
  signal lineLoader_wayToAllocate_willIncrement : std_logic;
  signal lineLoader_wayToAllocate_willClear : std_logic;
  signal lineLoader_wayToAllocate_willOverflowIfInc : std_logic;
  signal lineLoader_wayToAllocate_willOverflow : std_logic;
  signal lineLoader_wordIndex : unsigned(2 downto 0);
  attribute keep of lineLoader_wordIndex : signal is true;
  attribute syn_keep of lineLoader_wordIndex : signal is true;
  signal lineLoader_write_tag_0_valid : std_logic;
  signal lineLoader_write_tag_0_payload_address : unsigned(7 downto 0);
  signal lineLoader_write_tag_0_payload_data_valid : std_logic;
  signal lineLoader_write_tag_0_payload_data_error : std_logic;
  signal lineLoader_write_tag_0_payload_data_address : unsigned(18 downto 0);
  signal lineLoader_write_data_0_valid : std_logic;
  signal lineLoader_write_data_0_payload_address : unsigned(10 downto 0);
  signal lineLoader_write_data_0_payload_data : std_logic_vector(31 downto 0);
  signal when_InstructionCache_l401 : std_logic;
  signal zz_fetchStage_read_banksValue_0_dataMem : unsigned(10 downto 0);
  signal zz_fetchStage_read_banksValue_0_dataMem_1 : std_logic;
  signal fetchStage_read_banksValue_0_dataMem : std_logic_vector(31 downto 0);
  signal fetchStage_read_banksValue_0_data : std_logic_vector(31 downto 0);
  signal zz_fetchStage_read_waysValues_0_tag_valid : unsigned(7 downto 0);
  signal zz_fetchStage_read_waysValues_0_tag_valid_1 : std_logic;
  signal fetchStage_read_waysValues_0_tag_valid : std_logic;
  signal fetchStage_read_waysValues_0_tag_error : std_logic;
  signal fetchStage_read_waysValues_0_tag_address : unsigned(18 downto 0);
  signal zz_fetchStage_read_waysValues_0_tag_valid_2 : std_logic_vector(20 downto 0);
  signal fetchStage_hit_hits_0 : std_logic;
  signal fetchStage_hit_valid : std_logic;
  signal fetchStage_hit_error : std_logic;
  signal fetchStage_hit_data : std_logic_vector(31 downto 0);
  signal fetchStage_hit_word : std_logic_vector(31 downto 0);
  signal when_InstructionCache_l435 : std_logic;
  signal io_cpu_fetch_data_regNextWhen : std_logic_vector(31 downto 0);
  signal when_InstructionCache_l459 : std_logic;
  signal decodeStage_mmuRsp_physicalAddress : unsigned(31 downto 0);
  signal decodeStage_mmuRsp_isIoAccess : std_logic;
  signal decodeStage_mmuRsp_isPaging : std_logic;
  signal decodeStage_mmuRsp_allowRead : std_logic;
  signal decodeStage_mmuRsp_allowWrite : std_logic;
  signal decodeStage_mmuRsp_allowExecute : std_logic;
  signal decodeStage_mmuRsp_exception : std_logic;
  signal decodeStage_mmuRsp_refilling : std_logic;
  signal decodeStage_mmuRsp_bypassTranslation : std_logic;
  signal when_InstructionCache_l459_1 : std_logic;
  signal decodeStage_hit_valid : std_logic;
  signal when_InstructionCache_l459_2 : std_logic;
  signal decodeStage_hit_error : std_logic;
  signal when_Fetcher_l398 : std_logic;
  type banks_0_type is array (0 to 2047) of std_logic_vector(31 downto 0);
  signal banks_0 : banks_0_type;
  type ways_0_tags_type is array (0 to 255) of std_logic_vector(20 downto 0);
  signal ways_0_tags : ways_0_tags_type;
begin
  io_mem_cmd_valid <= io_mem_cmd_valid_read_buffer;
  io_cpu_fetch_data <= io_cpu_fetch_data_read_buffer;
  zz_ways_0_tags_port <= pkg_cat(std_logic_vector(lineLoader_write_tag_0_payload_data_address),pkg_cat(pkg_toStdLogicVector(lineLoader_write_tag_0_payload_data_error),pkg_toStdLogicVector(lineLoader_write_tag_0_payload_data_valid)));
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_1 = '1' then
        banks_0(to_integer(lineLoader_write_data_0_payload_address)) <= lineLoader_write_data_0_payload_data;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_fetchStage_read_banksValue_0_dataMem_1 = '1' then
        zz_banks_0_port0 <= banks_0(to_integer(zz_fetchStage_read_banksValue_0_dataMem));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_2 = '1' then
        ways_0_tags(to_integer(lineLoader_write_tag_0_payload_address)) <= zz_ways_0_tags_port;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_fetchStage_read_waysValues_0_tag_valid_1 = '1' then
        zz_ways_0_tags_port0 <= ways_0_tags(to_integer(zz_fetchStage_read_waysValues_0_tag_valid));
      end if;
    end if;
  end process;

  process(lineLoader_write_data_0_valid)
  begin
    zz_1 <= pkg_toStdLogic(false);
    if lineLoader_write_data_0_valid = '1' then
      zz_1 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(lineLoader_write_tag_0_valid)
  begin
    zz_2 <= pkg_toStdLogic(false);
    if lineLoader_write_tag_0_valid = '1' then
      zz_2 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_mem_rsp_valid,when_InstructionCache_l401)
  begin
    lineLoader_fire <= pkg_toStdLogic(false);
    if io_mem_rsp_valid = '1' then
      if when_InstructionCache_l401 = '1' then
        lineLoader_fire <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  process(lineLoader_valid,lineLoader_flushPending,when_InstructionCache_l338,when_InstructionCache_l342,io_flush)
  begin
    io_cpu_prefetch_haltIt <= (lineLoader_valid or lineLoader_flushPending);
    if when_InstructionCache_l338 = '1' then
      io_cpu_prefetch_haltIt <= pkg_toStdLogic(true);
    end if;
    if when_InstructionCache_l342 = '1' then
      io_cpu_prefetch_haltIt <= pkg_toStdLogic(true);
    end if;
    if io_flush = '1' then
      io_cpu_prefetch_haltIt <= pkg_toStdLogic(true);
    end if;
  end process;

  when_InstructionCache_l338 <= (not pkg_extract(lineLoader_flushCounter,8));
  when_InstructionCache_l342 <= (not zz_when_InstructionCache_l342);
  when_InstructionCache_l351 <= (lineLoader_flushPending and (not (lineLoader_valid or io_cpu_fetch_isValid)));
  io_mem_cmd_fire <= (io_mem_cmd_valid_read_buffer and io_mem_cmd_ready);
  io_mem_cmd_valid_read_buffer <= (lineLoader_valid and (not lineLoader_cmdSent));
  io_mem_cmd_payload_address <= unsigned(pkg_cat(std_logic_vector(pkg_extract(lineLoader_address,31,5)),std_logic_vector(pkg_unsigned("00000"))));
  io_mem_cmd_payload_size <= pkg_unsigned("101");
  when_Utils_l485 <= (not lineLoader_valid);
  process(when_Utils_l485)
  begin
    lineLoader_wayToAllocate_willIncrement <= pkg_toStdLogic(false);
    if when_Utils_l485 = '1' then
      lineLoader_wayToAllocate_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  lineLoader_wayToAllocate_willClear <= pkg_toStdLogic(false);
  lineLoader_wayToAllocate_willOverflowIfInc <= pkg_toStdLogic(true);
  lineLoader_wayToAllocate_willOverflow <= (lineLoader_wayToAllocate_willOverflowIfInc and lineLoader_wayToAllocate_willIncrement);
  lineLoader_write_tag_0_valid <= ((pkg_toStdLogic(true) and lineLoader_fire) or (not pkg_extract(lineLoader_flushCounter,8)));
  lineLoader_write_tag_0_payload_address <= pkg_mux(pkg_extract(lineLoader_flushCounter,8),pkg_extract(lineLoader_address,12,5),pkg_extract(lineLoader_flushCounter,7,0));
  lineLoader_write_tag_0_payload_data_valid <= pkg_extract(lineLoader_flushCounter,8);
  lineLoader_write_tag_0_payload_data_error <= (lineLoader_hadError or io_mem_rsp_payload_error);
  lineLoader_write_tag_0_payload_data_address <= pkg_extract(lineLoader_address,31,13);
  lineLoader_write_data_0_valid <= (io_mem_rsp_valid and pkg_toStdLogic(true));
  lineLoader_write_data_0_payload_address <= unsigned(pkg_cat(std_logic_vector(pkg_extract(lineLoader_address,12,5)),std_logic_vector(lineLoader_wordIndex)));
  lineLoader_write_data_0_payload_data <= io_mem_rsp_payload_data;
  when_InstructionCache_l401 <= pkg_toStdLogic(lineLoader_wordIndex = pkg_unsigned("111"));
  zz_fetchStage_read_banksValue_0_dataMem <= pkg_extract(io_cpu_prefetch_pc,12,2);
  zz_fetchStage_read_banksValue_0_dataMem_1 <= (not io_cpu_fetch_isStuck);
  fetchStage_read_banksValue_0_dataMem <= zz_banks_0_port0;
  fetchStage_read_banksValue_0_data <= pkg_extract(fetchStage_read_banksValue_0_dataMem,31,0);
  zz_fetchStage_read_waysValues_0_tag_valid <= pkg_extract(io_cpu_prefetch_pc,12,5);
  zz_fetchStage_read_waysValues_0_tag_valid_1 <= (not io_cpu_fetch_isStuck);
  zz_fetchStage_read_waysValues_0_tag_valid_2 <= zz_ways_0_tags_port0;
  fetchStage_read_waysValues_0_tag_valid <= pkg_extract(zz_fetchStage_read_waysValues_0_tag_valid_2,0);
  fetchStage_read_waysValues_0_tag_error <= pkg_extract(zz_fetchStage_read_waysValues_0_tag_valid_2,1);
  fetchStage_read_waysValues_0_tag_address <= unsigned(pkg_extract(zz_fetchStage_read_waysValues_0_tag_valid_2,20,2));
  fetchStage_hit_hits_0 <= (fetchStage_read_waysValues_0_tag_valid and pkg_toStdLogic(fetchStage_read_waysValues_0_tag_address = pkg_extract(io_cpu_fetch_mmuRsp_physicalAddress,31,13)));
  fetchStage_hit_valid <= pkg_toStdLogic(pkg_toStdLogicVector(fetchStage_hit_hits_0) /= pkg_stdLogicVector("0"));
  fetchStage_hit_error <= fetchStage_read_waysValues_0_tag_error;
  fetchStage_hit_data <= fetchStage_read_banksValue_0_data;
  fetchStage_hit_word <= fetchStage_hit_data;
  io_cpu_fetch_data_read_buffer <= fetchStage_hit_word;
  when_InstructionCache_l435 <= (not io_cpu_decode_isStuck);
  io_cpu_decode_data <= io_cpu_fetch_data_regNextWhen;
  io_cpu_fetch_physicalAddress <= io_cpu_fetch_mmuRsp_physicalAddress;
  when_InstructionCache_l459 <= (not io_cpu_decode_isStuck);
  when_InstructionCache_l459_1 <= (not io_cpu_decode_isStuck);
  when_InstructionCache_l459_2 <= (not io_cpu_decode_isStuck);
  io_cpu_decode_cacheMiss <= (not decodeStage_hit_valid);
  io_cpu_decode_error <= (decodeStage_hit_error or ((not decodeStage_mmuRsp_isPaging) and (decodeStage_mmuRsp_exception or (not decodeStage_mmuRsp_allowExecute))));
  io_cpu_decode_mmuRefilling <= decodeStage_mmuRsp_refilling;
  io_cpu_decode_mmuException <= (((not decodeStage_mmuRsp_refilling) and decodeStage_mmuRsp_isPaging) and (decodeStage_mmuRsp_exception or (not decodeStage_mmuRsp_allowExecute)));
  io_cpu_decode_physicalAddress <= decodeStage_mmuRsp_physicalAddress;
  when_Fetcher_l398 <= pkg_toStdLogic(zz_when_Fetcher_l398 /= pkg_unsigned("000"));
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      lineLoader_valid <= pkg_toStdLogic(false);
      lineLoader_hadError <= pkg_toStdLogic(false);
      lineLoader_flushPending <= pkg_toStdLogic(true);
      lineLoader_cmdSent <= pkg_toStdLogic(false);
      lineLoader_wordIndex <= pkg_unsigned("000");
    elsif rising_edge(io_mainClk) then
      if lineLoader_fire = '1' then
        lineLoader_valid <= pkg_toStdLogic(false);
      end if;
      if lineLoader_fire = '1' then
        lineLoader_hadError <= pkg_toStdLogic(false);
      end if;
      if io_cpu_fill_valid = '1' then
        lineLoader_valid <= pkg_toStdLogic(true);
      end if;
      if io_flush = '1' then
        lineLoader_flushPending <= pkg_toStdLogic(true);
      end if;
      if when_InstructionCache_l351 = '1' then
        lineLoader_flushPending <= pkg_toStdLogic(false);
      end if;
      if io_mem_cmd_fire = '1' then
        lineLoader_cmdSent <= pkg_toStdLogic(true);
      end if;
      if lineLoader_fire = '1' then
        lineLoader_cmdSent <= pkg_toStdLogic(false);
      end if;
      if io_mem_rsp_valid = '1' then
        lineLoader_wordIndex <= (lineLoader_wordIndex + pkg_unsigned("001"));
        if io_mem_rsp_payload_error = '1' then
          lineLoader_hadError <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_cpu_fill_valid = '1' then
        lineLoader_address <= io_cpu_fill_payload;
      end if;
      if when_InstructionCache_l338 = '1' then
        lineLoader_flushCounter <= (lineLoader_flushCounter + pkg_unsigned("000000001"));
      end if;
      zz_when_InstructionCache_l342 <= pkg_extract(lineLoader_flushCounter,8);
      if when_InstructionCache_l351 = '1' then
        lineLoader_flushCounter <= pkg_unsigned("000000000");
      end if;
      if when_InstructionCache_l435 = '1' then
        io_cpu_fetch_data_regNextWhen <= io_cpu_fetch_data_read_buffer;
      end if;
      if when_InstructionCache_l459 = '1' then
        decodeStage_mmuRsp_physicalAddress <= io_cpu_fetch_mmuRsp_physicalAddress;
        decodeStage_mmuRsp_isIoAccess <= io_cpu_fetch_mmuRsp_isIoAccess;
        decodeStage_mmuRsp_isPaging <= io_cpu_fetch_mmuRsp_isPaging;
        decodeStage_mmuRsp_allowRead <= io_cpu_fetch_mmuRsp_allowRead;
        decodeStage_mmuRsp_allowWrite <= io_cpu_fetch_mmuRsp_allowWrite;
        decodeStage_mmuRsp_allowExecute <= io_cpu_fetch_mmuRsp_allowExecute;
        decodeStage_mmuRsp_exception <= io_cpu_fetch_mmuRsp_exception;
        decodeStage_mmuRsp_refilling <= io_cpu_fetch_mmuRsp_refilling;
        decodeStage_mmuRsp_bypassTranslation <= io_cpu_fetch_mmuRsp_bypassTranslation;
      end if;
      if when_InstructionCache_l459_1 = '1' then
        decodeStage_hit_valid <= fetchStage_hit_valid;
      end if;
      if when_InstructionCache_l459_2 = '1' then
        decodeStage_hit_error <= fetchStage_hit_error;
      end if;
      if when_Fetcher_l398 = '1' then
        io_cpu_fetch_data_regNextWhen <= zz_io_cpu_fetch_data_regNextWhen;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity DataCache is
  port(
    io_cpu_execute_isValid : in std_logic;
    io_cpu_execute_address : in unsigned(31 downto 0);
    io_cpu_execute_haltIt : out std_logic;
    io_cpu_execute_args_wr : in std_logic;
    io_cpu_execute_args_size : in unsigned(1 downto 0);
    io_cpu_execute_args_totalyConsistent : in std_logic;
    io_cpu_execute_refilling : out std_logic;
    io_cpu_memory_isValid : in std_logic;
    io_cpu_memory_isStuck : in std_logic;
    io_cpu_memory_isWrite : out std_logic;
    io_cpu_memory_address : in unsigned(31 downto 0);
    io_cpu_memory_mmuRsp_physicalAddress : in unsigned(31 downto 0);
    io_cpu_memory_mmuRsp_isIoAccess : in std_logic;
    io_cpu_memory_mmuRsp_isPaging : in std_logic;
    io_cpu_memory_mmuRsp_allowRead : in std_logic;
    io_cpu_memory_mmuRsp_allowWrite : in std_logic;
    io_cpu_memory_mmuRsp_allowExecute : in std_logic;
    io_cpu_memory_mmuRsp_exception : in std_logic;
    io_cpu_memory_mmuRsp_refilling : in std_logic;
    io_cpu_memory_mmuRsp_bypassTranslation : in std_logic;
    io_cpu_writeBack_isValid : in std_logic;
    io_cpu_writeBack_isStuck : in std_logic;
    io_cpu_writeBack_isUser : in std_logic;
    io_cpu_writeBack_haltIt : out std_logic;
    io_cpu_writeBack_isWrite : out std_logic;
    io_cpu_writeBack_storeData : in std_logic_vector(31 downto 0);
    io_cpu_writeBack_data : out std_logic_vector(31 downto 0);
    io_cpu_writeBack_address : in unsigned(31 downto 0);
    io_cpu_writeBack_mmuException : out std_logic;
    io_cpu_writeBack_unalignedAccess : out std_logic;
    io_cpu_writeBack_accessError : out std_logic;
    io_cpu_writeBack_keepMemRspData : out std_logic;
    io_cpu_writeBack_fence_SW : in std_logic;
    io_cpu_writeBack_fence_SR : in std_logic;
    io_cpu_writeBack_fence_SO : in std_logic;
    io_cpu_writeBack_fence_SI : in std_logic;
    io_cpu_writeBack_fence_PW : in std_logic;
    io_cpu_writeBack_fence_PR : in std_logic;
    io_cpu_writeBack_fence_PO : in std_logic;
    io_cpu_writeBack_fence_PI : in std_logic;
    io_cpu_writeBack_fence_FM : in std_logic_vector(3 downto 0);
    io_cpu_writeBack_exclusiveOk : out std_logic;
    io_cpu_redo : out std_logic;
    io_cpu_flush_valid : in std_logic;
    io_cpu_flush_ready : out std_logic;
    io_mem_cmd_valid : out std_logic;
    io_mem_cmd_ready : in std_logic;
    io_mem_cmd_payload_wr : out std_logic;
    io_mem_cmd_payload_uncached : out std_logic;
    io_mem_cmd_payload_address : out unsigned(31 downto 0);
    io_mem_cmd_payload_data : out std_logic_vector(31 downto 0);
    io_mem_cmd_payload_mask : out std_logic_vector(3 downto 0);
    io_mem_cmd_payload_size : out unsigned(2 downto 0);
    io_mem_cmd_payload_last : out std_logic;
    io_mem_rsp_valid : in std_logic;
    io_mem_rsp_payload_last : in std_logic;
    io_mem_rsp_payload_data : in std_logic_vector(31 downto 0);
    io_mem_rsp_payload_error : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end DataCache;

architecture arch of DataCache is
  signal zz_ways_0_tags_port0 : std_logic_vector(22 downto 0);
  signal zz_ways_0_data_port0 : std_logic_vector(31 downto 0);
  signal zz_ways_1_tags_port0 : std_logic_vector(22 downto 0);
  signal zz_ways_1_data_port0 : std_logic_vector(31 downto 0);
  signal zz_ways_2_tags_port0 : std_logic_vector(22 downto 0);
  signal zz_ways_2_data_port0 : std_logic_vector(31 downto 0);
  signal zz_ways_3_tags_port0 : std_logic_vector(22 downto 0);
  signal zz_ways_3_data_port0 : std_logic_vector(31 downto 0);
  signal io_mem_cmd_valid_read_buffer : std_logic;
  signal io_cpu_flush_ready_read_buffer : std_logic;
  signal io_cpu_redo_read_buffer : std_logic;
  signal io_cpu_writeBack_accessError_read_buffer : std_logic;
  signal io_cpu_writeBack_mmuException_read_buffer : std_logic;
  signal io_cpu_writeBack_unalignedAccess_read_buffer : std_logic;
  signal io_cpu_writeBack_haltIt_read_buffer : std_logic;
  signal zz_ways_0_tags_port : std_logic_vector(22 downto 0);
  signal zz_ways_1_tags_port : std_logic_vector(22 downto 0);
  signal zz_ways_2_tags_port : std_logic_vector(22 downto 0);
  signal zz_ways_3_tags_port : std_logic_vector(22 downto 0);
  signal zz_stageB_dataMux_3 : std_logic_vector(31 downto 0);
  signal zz_stageB_dataMux_4 : unsigned(1 downto 0);

  signal zz_1 : std_logic;
  signal zz_2 : std_logic;
  signal zz_3 : std_logic;
  signal zz_4 : std_logic;
  signal zz_5 : std_logic;
  signal zz_6 : std_logic;
  signal zz_7 : std_logic;
  signal zz_8 : std_logic;
  signal haltCpu : std_logic;
  signal tagsReadCmd_valid : std_logic;
  signal tagsReadCmd_payload : unsigned(5 downto 0);
  signal tagsWriteCmd_valid : std_logic;
  signal tagsWriteCmd_payload_way : std_logic_vector(3 downto 0);
  signal tagsWriteCmd_payload_address : unsigned(5 downto 0);
  signal tagsWriteCmd_payload_data_valid : std_logic;
  signal tagsWriteCmd_payload_data_error : std_logic;
  signal tagsWriteCmd_payload_data_address : unsigned(20 downto 0);
  signal tagsWriteLastCmd_valid : std_logic;
  signal tagsWriteLastCmd_payload_way : std_logic_vector(3 downto 0);
  signal tagsWriteLastCmd_payload_address : unsigned(5 downto 0);
  signal tagsWriteLastCmd_payload_data_valid : std_logic;
  signal tagsWriteLastCmd_payload_data_error : std_logic;
  signal tagsWriteLastCmd_payload_data_address : unsigned(20 downto 0);
  signal dataReadCmd_valid : std_logic;
  signal dataReadCmd_payload : unsigned(8 downto 0);
  signal dataWriteCmd_valid : std_logic;
  signal dataWriteCmd_payload_way : std_logic_vector(3 downto 0);
  signal dataWriteCmd_payload_address : unsigned(8 downto 0);
  signal dataWriteCmd_payload_data : std_logic_vector(31 downto 0);
  signal dataWriteCmd_payload_mask : std_logic_vector(3 downto 0);
  signal zz_ways_0_tagsReadRsp_valid : std_logic;
  signal ways_0_tagsReadRsp_valid : std_logic;
  signal ways_0_tagsReadRsp_error : std_logic;
  signal ways_0_tagsReadRsp_address : unsigned(20 downto 0);
  signal zz_ways_0_tagsReadRsp_valid_1 : std_logic_vector(22 downto 0);
  signal zz_ways_0_dataReadRspMem : std_logic;
  signal ways_0_dataReadRspMem : std_logic_vector(31 downto 0);
  signal ways_0_dataReadRsp : std_logic_vector(31 downto 0);
  signal when_DataCache_l635 : std_logic;
  signal when_DataCache_l638 : std_logic;
  signal zz_ways_1_tagsReadRsp_valid : std_logic;
  signal ways_1_tagsReadRsp_valid : std_logic;
  signal ways_1_tagsReadRsp_error : std_logic;
  signal ways_1_tagsReadRsp_address : unsigned(20 downto 0);
  signal zz_ways_1_tagsReadRsp_valid_1 : std_logic_vector(22 downto 0);
  signal zz_ways_1_dataReadRspMem : std_logic;
  signal ways_1_dataReadRspMem : std_logic_vector(31 downto 0);
  signal ways_1_dataReadRsp : std_logic_vector(31 downto 0);
  signal when_DataCache_l635_1 : std_logic;
  signal when_DataCache_l638_1 : std_logic;
  signal zz_ways_2_tagsReadRsp_valid : std_logic;
  signal ways_2_tagsReadRsp_valid : std_logic;
  signal ways_2_tagsReadRsp_error : std_logic;
  signal ways_2_tagsReadRsp_address : unsigned(20 downto 0);
  signal zz_ways_2_tagsReadRsp_valid_1 : std_logic_vector(22 downto 0);
  signal zz_ways_2_dataReadRspMem : std_logic;
  signal ways_2_dataReadRspMem : std_logic_vector(31 downto 0);
  signal ways_2_dataReadRsp : std_logic_vector(31 downto 0);
  signal when_DataCache_l635_2 : std_logic;
  signal when_DataCache_l638_2 : std_logic;
  signal zz_ways_3_tagsReadRsp_valid : std_logic;
  signal ways_3_tagsReadRsp_valid : std_logic;
  signal ways_3_tagsReadRsp_error : std_logic;
  signal ways_3_tagsReadRsp_address : unsigned(20 downto 0);
  signal zz_ways_3_tagsReadRsp_valid_1 : std_logic_vector(22 downto 0);
  signal zz_ways_3_dataReadRspMem : std_logic;
  signal ways_3_dataReadRspMem : std_logic_vector(31 downto 0);
  signal ways_3_dataReadRsp : std_logic_vector(31 downto 0);
  signal when_DataCache_l635_3 : std_logic;
  signal when_DataCache_l638_3 : std_logic;
  signal when_DataCache_l657 : std_logic;
  signal rspSync : std_logic;
  signal rspLast : std_logic;
  signal memCmdSent : std_logic;
  signal io_mem_cmd_fire : std_logic;
  signal when_DataCache_l679 : std_logic;
  signal zz_stage0_mask : std_logic_vector(3 downto 0);
  signal stage0_mask : std_logic_vector(3 downto 0);
  signal stage0_dataColisions : std_logic_vector(3 downto 0);
  signal zz_stage0_dataColisions : unsigned(8 downto 0);
  signal zz_stage0_dataColisions_1 : std_logic_vector(3 downto 0);
  signal stage0_wayInvalidate : std_logic_vector(3 downto 0);
  signal stage0_isAmo : std_logic;
  signal when_DataCache_l764 : std_logic;
  signal stageA_request_wr : std_logic;
  signal stageA_request_size : unsigned(1 downto 0);
  signal stageA_request_totalyConsistent : std_logic;
  signal when_DataCache_l764_1 : std_logic;
  signal stageA_mask : std_logic_vector(3 downto 0);
  signal stageA_isAmo : std_logic;
  signal stageA_isLrsc : std_logic;
  signal stageA_wayHits : std_logic_vector(3 downto 0);
  signal when_DataCache_l764_2 : std_logic;
  signal stageA_wayInvalidate : std_logic_vector(3 downto 0);
  signal when_DataCache_l764_3 : std_logic;
  signal stage0_dataColisions_regNextWhen : std_logic_vector(3 downto 0);
  signal zz_stageA_dataColisions : std_logic_vector(3 downto 0);
  signal zz_stageA_dataColisions_1 : unsigned(8 downto 0);
  signal zz_stageA_dataColisions_2 : std_logic_vector(3 downto 0);
  signal stageA_dataColisions : std_logic_vector(3 downto 0);
  signal when_DataCache_l815 : std_logic;
  signal stageB_request_wr : std_logic;
  signal stageB_request_size : unsigned(1 downto 0);
  signal stageB_request_totalyConsistent : std_logic;
  signal stageB_mmuRspFreeze : std_logic;
  signal when_DataCache_l817 : std_logic;
  signal stageB_mmuRsp_physicalAddress : unsigned(31 downto 0);
  signal stageB_mmuRsp_isIoAccess : std_logic;
  signal stageB_mmuRsp_isPaging : std_logic;
  signal stageB_mmuRsp_allowRead : std_logic;
  signal stageB_mmuRsp_allowWrite : std_logic;
  signal stageB_mmuRsp_allowExecute : std_logic;
  signal stageB_mmuRsp_exception : std_logic;
  signal stageB_mmuRsp_refilling : std_logic;
  signal stageB_mmuRsp_bypassTranslation : std_logic;
  signal when_DataCache_l814 : std_logic;
  signal stageB_tagsReadRsp_0_valid : std_logic;
  signal stageB_tagsReadRsp_0_error : std_logic;
  signal stageB_tagsReadRsp_0_address : unsigned(20 downto 0);
  signal when_DataCache_l814_1 : std_logic;
  signal stageB_tagsReadRsp_1_valid : std_logic;
  signal stageB_tagsReadRsp_1_error : std_logic;
  signal stageB_tagsReadRsp_1_address : unsigned(20 downto 0);
  signal when_DataCache_l814_2 : std_logic;
  signal stageB_tagsReadRsp_2_valid : std_logic;
  signal stageB_tagsReadRsp_2_error : std_logic;
  signal stageB_tagsReadRsp_2_address : unsigned(20 downto 0);
  signal when_DataCache_l814_3 : std_logic;
  signal stageB_tagsReadRsp_3_valid : std_logic;
  signal stageB_tagsReadRsp_3_error : std_logic;
  signal stageB_tagsReadRsp_3_address : unsigned(20 downto 0);
  signal when_DataCache_l814_4 : std_logic;
  signal stageB_dataReadRsp_0 : std_logic_vector(31 downto 0);
  signal when_DataCache_l814_5 : std_logic;
  signal stageB_dataReadRsp_1 : std_logic_vector(31 downto 0);
  signal when_DataCache_l814_6 : std_logic;
  signal stageB_dataReadRsp_2 : std_logic_vector(31 downto 0);
  signal when_DataCache_l814_7 : std_logic;
  signal stageB_dataReadRsp_3 : std_logic_vector(31 downto 0);
  signal when_DataCache_l813 : std_logic;
  signal stageB_wayInvalidate : std_logic_vector(3 downto 0);
  signal stageB_consistancyHazard : std_logic;
  signal when_DataCache_l813_1 : std_logic;
  signal stageB_dataColisions : std_logic_vector(3 downto 0);
  signal when_DataCache_l813_2 : std_logic;
  signal stageB_unaligned : std_logic;
  signal when_DataCache_l813_3 : std_logic;
  signal stageB_waysHitsBeforeInvalidate : std_logic_vector(3 downto 0);
  signal stageB_waysHits : std_logic_vector(3 downto 0);
  signal stageB_waysHit : std_logic;
  signal zz_stageB_dataMux : std_logic;
  signal zz_stageB_dataMux_1 : std_logic;
  signal zz_stageB_dataMux_2 : std_logic;
  signal stageB_dataMux : std_logic_vector(31 downto 0);
  signal when_DataCache_l813_4 : std_logic;
  signal stageB_mask : std_logic_vector(3 downto 0);
  signal stageB_loaderValid : std_logic;
  signal stageB_ioMemRspMuxed : std_logic_vector(31 downto 0);
  signal stageB_flusher_waitDone : std_logic;
  signal stageB_flusher_hold : std_logic;
  signal stageB_flusher_counter : unsigned(6 downto 0);
  signal when_DataCache_l843 : std_logic;
  signal when_DataCache_l849 : std_logic;
  signal stageB_flusher_start : std_logic;
  signal stageB_isAmo : std_logic;
  signal stageB_isAmoCached : std_logic;
  signal stageB_isExternalLsrc : std_logic;
  signal stageB_isExternalAmo : std_logic;
  signal stageB_requestDataBypass : std_logic_vector(31 downto 0);
  signal stageB_cpuWriteToCache : std_logic;
  signal when_DataCache_l912 : std_logic;
  signal stageB_badPermissions : std_logic;
  signal stageB_loadStoreFault : std_logic;
  signal stageB_bypassCache : std_logic;
  signal when_DataCache_l981 : std_logic;
  signal when_DataCache_l990 : std_logic;
  signal when_DataCache_l995 : std_logic;
  signal when_DataCache_l1006 : std_logic;
  signal when_DataCache_l1018 : std_logic;
  signal when_DataCache_l977 : std_logic;
  signal when_DataCache_l1052 : std_logic;
  signal when_DataCache_l1061 : std_logic;
  signal loader_valid : std_logic;
  signal loader_counter_willIncrement : std_logic;
  signal loader_counter_willClear : std_logic;
  signal loader_counter_valueNext : unsigned(2 downto 0);
  signal loader_counter_value : unsigned(2 downto 0);
  signal loader_counter_willOverflowIfInc : std_logic;
  signal loader_counter_willOverflow : std_logic;
  signal loader_waysAllocator : std_logic_vector(3 downto 0);
  signal loader_error : std_logic;
  signal loader_kill : std_logic;
  signal loader_killReg : std_logic;
  signal when_DataCache_l1076 : std_logic;
  signal loader_done : std_logic;
  signal when_DataCache_l1104 : std_logic;
  signal loader_valid_regNext : std_logic;
  signal when_DataCache_l1108 : std_logic;
  signal when_DataCache_l1111 : std_logic;
  type ways_0_tags_type is array (0 to 63) of std_logic_vector(22 downto 0);
  signal ways_0_tags : ways_0_tags_type;
  type ways_0_data_type is array (0 to 511) of std_logic_vector(7 downto 0);
  signal ways_0_data_symbol0 : ways_0_data_type;
  signal ways_0_data_symbol1 : ways_0_data_type;
  signal ways_0_data_symbol2 : ways_0_data_type;
  signal ways_0_data_symbol3 : ways_0_data_type;
  signal zz_9 : std_logic_vector(7 downto 0);
  signal zz_10 : std_logic_vector(7 downto 0);
  signal zz_11 : std_logic_vector(7 downto 0);
  signal zz_12 : std_logic_vector(7 downto 0);
  type ways_1_tags_type is array (0 to 63) of std_logic_vector(22 downto 0);
  signal ways_1_tags : ways_1_tags_type;
  type ways_1_data_type is array (0 to 511) of std_logic_vector(7 downto 0);
  signal ways_1_data_symbol0 : ways_1_data_type;
  signal ways_1_data_symbol1 : ways_1_data_type;
  signal ways_1_data_symbol2 : ways_1_data_type;
  signal ways_1_data_symbol3 : ways_1_data_type;
  signal zz_13 : std_logic_vector(7 downto 0);
  signal zz_14 : std_logic_vector(7 downto 0);
  signal zz_15 : std_logic_vector(7 downto 0);
  signal zz_16 : std_logic_vector(7 downto 0);
  type ways_2_tags_type is array (0 to 63) of std_logic_vector(22 downto 0);
  signal ways_2_tags : ways_2_tags_type;
  type ways_2_data_type is array (0 to 511) of std_logic_vector(7 downto 0);
  signal ways_2_data_symbol0 : ways_2_data_type;
  signal ways_2_data_symbol1 : ways_2_data_type;
  signal ways_2_data_symbol2 : ways_2_data_type;
  signal ways_2_data_symbol3 : ways_2_data_type;
  signal zz_17 : std_logic_vector(7 downto 0);
  signal zz_18 : std_logic_vector(7 downto 0);
  signal zz_19 : std_logic_vector(7 downto 0);
  signal zz_20 : std_logic_vector(7 downto 0);
  type ways_3_tags_type is array (0 to 63) of std_logic_vector(22 downto 0);
  signal ways_3_tags : ways_3_tags_type;
  type ways_3_data_type is array (0 to 511) of std_logic_vector(7 downto 0);
  signal ways_3_data_symbol0 : ways_3_data_type;
  signal ways_3_data_symbol1 : ways_3_data_type;
  signal ways_3_data_symbol2 : ways_3_data_type;
  signal ways_3_data_symbol3 : ways_3_data_type;
  signal zz_21 : std_logic_vector(7 downto 0);
  signal zz_22 : std_logic_vector(7 downto 0);
  signal zz_23 : std_logic_vector(7 downto 0);
  signal zz_24 : std_logic_vector(7 downto 0);
begin
  io_mem_cmd_valid <= io_mem_cmd_valid_read_buffer;
  io_cpu_flush_ready <= io_cpu_flush_ready_read_buffer;
  io_cpu_redo <= io_cpu_redo_read_buffer;
  io_cpu_writeBack_accessError <= io_cpu_writeBack_accessError_read_buffer;
  io_cpu_writeBack_mmuException <= io_cpu_writeBack_mmuException_read_buffer;
  io_cpu_writeBack_unalignedAccess <= io_cpu_writeBack_unalignedAccess_read_buffer;
  io_cpu_writeBack_haltIt <= io_cpu_writeBack_haltIt_read_buffer;
  zz_ways_0_tags_port <= pkg_cat(std_logic_vector(tagsWriteCmd_payload_data_address),pkg_cat(pkg_toStdLogicVector(tagsWriteCmd_payload_data_error),pkg_toStdLogicVector(tagsWriteCmd_payload_data_valid)));
  zz_ways_1_tags_port <= pkg_cat(std_logic_vector(tagsWriteCmd_payload_data_address),pkg_cat(pkg_toStdLogicVector(tagsWriteCmd_payload_data_error),pkg_toStdLogicVector(tagsWriteCmd_payload_data_valid)));
  zz_ways_2_tags_port <= pkg_cat(std_logic_vector(tagsWriteCmd_payload_data_address),pkg_cat(pkg_toStdLogicVector(tagsWriteCmd_payload_data_error),pkg_toStdLogicVector(tagsWriteCmd_payload_data_valid)));
  zz_ways_3_tags_port <= pkg_cat(std_logic_vector(tagsWriteCmd_payload_data_address),pkg_cat(pkg_toStdLogicVector(tagsWriteCmd_payload_data_error),pkg_toStdLogicVector(tagsWriteCmd_payload_data_valid)));
  zz_stageB_dataMux_4 <= unsigned(pkg_cat(pkg_toStdLogicVector(zz_stageB_dataMux_2),pkg_toStdLogicVector(zz_stageB_dataMux_1)));
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_0_tagsReadRsp_valid = '1' then
        zz_ways_0_tags_port0 <= ways_0_tags(to_integer(tagsReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_8 = '1' then
        ways_0_tags(to_integer(tagsWriteCmd_payload_address)) <= zz_ways_0_tags_port;
      end if;
    end if;
  end process;

  process (zz_9, zz_10, zz_11, zz_12)
  begin
    zz_ways_0_data_port0 <= zz_12 & zz_11 & zz_10 & zz_9;
  end process;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_0_dataReadRspMem = '1' then
        zz_9 <= ways_0_data_symbol0(to_integer(dataReadCmd_payload));
        zz_10 <= ways_0_data_symbol1(to_integer(dataReadCmd_payload));
        zz_11 <= ways_0_data_symbol2(to_integer(dataReadCmd_payload));
        zz_12 <= ways_0_data_symbol3(to_integer(dataReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if dataWriteCmd_payload_mask(0) = '1' and zz_7 = '1' then
        ways_0_data_symbol0(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(7 downto 0);
      end if;
      if dataWriteCmd_payload_mask(1) = '1' and zz_7 = '1' then
        ways_0_data_symbol1(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(15 downto 8);
      end if;
      if dataWriteCmd_payload_mask(2) = '1' and zz_7 = '1' then
        ways_0_data_symbol2(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(23 downto 16);
      end if;
      if dataWriteCmd_payload_mask(3) = '1' and zz_7 = '1' then
        ways_0_data_symbol3(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(31 downto 24);
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_1_tagsReadRsp_valid = '1' then
        zz_ways_1_tags_port0 <= ways_1_tags(to_integer(tagsReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_6 = '1' then
        ways_1_tags(to_integer(tagsWriteCmd_payload_address)) <= zz_ways_1_tags_port;
      end if;
    end if;
  end process;

  process (zz_13, zz_14, zz_15, zz_16)
  begin
    zz_ways_1_data_port0 <= zz_16 & zz_15 & zz_14 & zz_13;
  end process;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_1_dataReadRspMem = '1' then
        zz_13 <= ways_1_data_symbol0(to_integer(dataReadCmd_payload));
        zz_14 <= ways_1_data_symbol1(to_integer(dataReadCmd_payload));
        zz_15 <= ways_1_data_symbol2(to_integer(dataReadCmd_payload));
        zz_16 <= ways_1_data_symbol3(to_integer(dataReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if dataWriteCmd_payload_mask(0) = '1' and zz_5 = '1' then
        ways_1_data_symbol0(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(7 downto 0);
      end if;
      if dataWriteCmd_payload_mask(1) = '1' and zz_5 = '1' then
        ways_1_data_symbol1(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(15 downto 8);
      end if;
      if dataWriteCmd_payload_mask(2) = '1' and zz_5 = '1' then
        ways_1_data_symbol2(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(23 downto 16);
      end if;
      if dataWriteCmd_payload_mask(3) = '1' and zz_5 = '1' then
        ways_1_data_symbol3(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(31 downto 24);
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_2_tagsReadRsp_valid = '1' then
        zz_ways_2_tags_port0 <= ways_2_tags(to_integer(tagsReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_4 = '1' then
        ways_2_tags(to_integer(tagsWriteCmd_payload_address)) <= zz_ways_2_tags_port;
      end if;
    end if;
  end process;

  process (zz_17, zz_18, zz_19, zz_20)
  begin
    zz_ways_2_data_port0 <= zz_20 & zz_19 & zz_18 & zz_17;
  end process;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_2_dataReadRspMem = '1' then
        zz_17 <= ways_2_data_symbol0(to_integer(dataReadCmd_payload));
        zz_18 <= ways_2_data_symbol1(to_integer(dataReadCmd_payload));
        zz_19 <= ways_2_data_symbol2(to_integer(dataReadCmd_payload));
        zz_20 <= ways_2_data_symbol3(to_integer(dataReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if dataWriteCmd_payload_mask(0) = '1' and zz_3 = '1' then
        ways_2_data_symbol0(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(7 downto 0);
      end if;
      if dataWriteCmd_payload_mask(1) = '1' and zz_3 = '1' then
        ways_2_data_symbol1(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(15 downto 8);
      end if;
      if dataWriteCmd_payload_mask(2) = '1' and zz_3 = '1' then
        ways_2_data_symbol2(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(23 downto 16);
      end if;
      if dataWriteCmd_payload_mask(3) = '1' and zz_3 = '1' then
        ways_2_data_symbol3(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(31 downto 24);
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_3_tagsReadRsp_valid = '1' then
        zz_ways_3_tags_port0 <= ways_3_tags(to_integer(tagsReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_2 = '1' then
        ways_3_tags(to_integer(tagsWriteCmd_payload_address)) <= zz_ways_3_tags_port;
      end if;
    end if;
  end process;

  process (zz_21, zz_22, zz_23, zz_24)
  begin
    zz_ways_3_data_port0 <= zz_24 & zz_23 & zz_22 & zz_21;
  end process;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_ways_3_dataReadRspMem = '1' then
        zz_21 <= ways_3_data_symbol0(to_integer(dataReadCmd_payload));
        zz_22 <= ways_3_data_symbol1(to_integer(dataReadCmd_payload));
        zz_23 <= ways_3_data_symbol2(to_integer(dataReadCmd_payload));
        zz_24 <= ways_3_data_symbol3(to_integer(dataReadCmd_payload));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if dataWriteCmd_payload_mask(0) = '1' and zz_1 = '1' then
        ways_3_data_symbol0(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(7 downto 0);
      end if;
      if dataWriteCmd_payload_mask(1) = '1' and zz_1 = '1' then
        ways_3_data_symbol1(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(15 downto 8);
      end if;
      if dataWriteCmd_payload_mask(2) = '1' and zz_1 = '1' then
        ways_3_data_symbol2(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(23 downto 16);
      end if;
      if dataWriteCmd_payload_mask(3) = '1' and zz_1 = '1' then
        ways_3_data_symbol3(to_integer(dataWriteCmd_payload_address)) <= dataWriteCmd_payload_data(31 downto 24);
      end if;
    end if;
  end process;

  process(zz_stageB_dataMux_4,stageB_dataReadRsp_0,stageB_dataReadRsp_1,stageB_dataReadRsp_2,stageB_dataReadRsp_3)
  begin
    case zz_stageB_dataMux_4 is
      when "00" =>
        zz_stageB_dataMux_3 <= stageB_dataReadRsp_0;
      when "01" =>
        zz_stageB_dataMux_3 <= stageB_dataReadRsp_1;
      when "10" =>
        zz_stageB_dataMux_3 <= stageB_dataReadRsp_2;
      when others =>
        zz_stageB_dataMux_3 <= stageB_dataReadRsp_3;
    end case;
  end process;

  process(when_DataCache_l638_3)
  begin
    zz_1 <= pkg_toStdLogic(false);
    if when_DataCache_l638_3 = '1' then
      zz_1 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l635_3)
  begin
    zz_2 <= pkg_toStdLogic(false);
    if when_DataCache_l635_3 = '1' then
      zz_2 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l638_2)
  begin
    zz_3 <= pkg_toStdLogic(false);
    if when_DataCache_l638_2 = '1' then
      zz_3 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l635_2)
  begin
    zz_4 <= pkg_toStdLogic(false);
    if when_DataCache_l635_2 = '1' then
      zz_4 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l638_1)
  begin
    zz_5 <= pkg_toStdLogic(false);
    if when_DataCache_l638_1 = '1' then
      zz_5 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l635_1)
  begin
    zz_6 <= pkg_toStdLogic(false);
    if when_DataCache_l635_1 = '1' then
      zz_6 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l638)
  begin
    zz_7 <= pkg_toStdLogic(false);
    if when_DataCache_l638 = '1' then
      zz_7 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l635)
  begin
    zz_8 <= pkg_toStdLogic(false);
    if when_DataCache_l635 = '1' then
      zz_8 <= pkg_toStdLogic(true);
    end if;
  end process;

  haltCpu <= pkg_toStdLogic(false);
  zz_ways_0_tagsReadRsp_valid <= (tagsReadCmd_valid and (not io_cpu_memory_isStuck));
  zz_ways_0_tagsReadRsp_valid_1 <= zz_ways_0_tags_port0;
  ways_0_tagsReadRsp_valid <= pkg_extract(zz_ways_0_tagsReadRsp_valid_1,0);
  ways_0_tagsReadRsp_error <= pkg_extract(zz_ways_0_tagsReadRsp_valid_1,1);
  ways_0_tagsReadRsp_address <= unsigned(pkg_extract(zz_ways_0_tagsReadRsp_valid_1,22,2));
  zz_ways_0_dataReadRspMem <= (dataReadCmd_valid and (not io_cpu_memory_isStuck));
  ways_0_dataReadRspMem <= zz_ways_0_data_port0;
  ways_0_dataReadRsp <= pkg_extract(ways_0_dataReadRspMem,31,0);
  when_DataCache_l635 <= (tagsWriteCmd_valid and pkg_extract(tagsWriteCmd_payload_way,0));
  when_DataCache_l638 <= (dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,0));
  zz_ways_1_tagsReadRsp_valid <= (tagsReadCmd_valid and (not io_cpu_memory_isStuck));
  zz_ways_1_tagsReadRsp_valid_1 <= zz_ways_1_tags_port0;
  ways_1_tagsReadRsp_valid <= pkg_extract(zz_ways_1_tagsReadRsp_valid_1,0);
  ways_1_tagsReadRsp_error <= pkg_extract(zz_ways_1_tagsReadRsp_valid_1,1);
  ways_1_tagsReadRsp_address <= unsigned(pkg_extract(zz_ways_1_tagsReadRsp_valid_1,22,2));
  zz_ways_1_dataReadRspMem <= (dataReadCmd_valid and (not io_cpu_memory_isStuck));
  ways_1_dataReadRspMem <= zz_ways_1_data_port0;
  ways_1_dataReadRsp <= pkg_extract(ways_1_dataReadRspMem,31,0);
  when_DataCache_l635_1 <= (tagsWriteCmd_valid and pkg_extract(tagsWriteCmd_payload_way,1));
  when_DataCache_l638_1 <= (dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,1));
  zz_ways_2_tagsReadRsp_valid <= (tagsReadCmd_valid and (not io_cpu_memory_isStuck));
  zz_ways_2_tagsReadRsp_valid_1 <= zz_ways_2_tags_port0;
  ways_2_tagsReadRsp_valid <= pkg_extract(zz_ways_2_tagsReadRsp_valid_1,0);
  ways_2_tagsReadRsp_error <= pkg_extract(zz_ways_2_tagsReadRsp_valid_1,1);
  ways_2_tagsReadRsp_address <= unsigned(pkg_extract(zz_ways_2_tagsReadRsp_valid_1,22,2));
  zz_ways_2_dataReadRspMem <= (dataReadCmd_valid and (not io_cpu_memory_isStuck));
  ways_2_dataReadRspMem <= zz_ways_2_data_port0;
  ways_2_dataReadRsp <= pkg_extract(ways_2_dataReadRspMem,31,0);
  when_DataCache_l635_2 <= (tagsWriteCmd_valid and pkg_extract(tagsWriteCmd_payload_way,2));
  when_DataCache_l638_2 <= (dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,2));
  zz_ways_3_tagsReadRsp_valid <= (tagsReadCmd_valid and (not io_cpu_memory_isStuck));
  zz_ways_3_tagsReadRsp_valid_1 <= zz_ways_3_tags_port0;
  ways_3_tagsReadRsp_valid <= pkg_extract(zz_ways_3_tagsReadRsp_valid_1,0);
  ways_3_tagsReadRsp_error <= pkg_extract(zz_ways_3_tagsReadRsp_valid_1,1);
  ways_3_tagsReadRsp_address <= unsigned(pkg_extract(zz_ways_3_tagsReadRsp_valid_1,22,2));
  zz_ways_3_dataReadRspMem <= (dataReadCmd_valid and (not io_cpu_memory_isStuck));
  ways_3_dataReadRspMem <= zz_ways_3_data_port0;
  ways_3_dataReadRsp <= pkg_extract(ways_3_dataReadRspMem,31,0);
  when_DataCache_l635_3 <= (tagsWriteCmd_valid and pkg_extract(tagsWriteCmd_payload_way,3));
  when_DataCache_l638_3 <= (dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,3));
  process(when_DataCache_l657)
  begin
    tagsReadCmd_valid <= pkg_toStdLogic(false);
    if when_DataCache_l657 = '1' then
      tagsReadCmd_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l657,io_cpu_execute_address)
  begin
    tagsReadCmd_payload <= pkg_unsigned("XXXXXX");
    if when_DataCache_l657 = '1' then
      tagsReadCmd_payload <= pkg_extract(io_cpu_execute_address,10,5);
    end if;
  end process;

  process(when_DataCache_l657)
  begin
    dataReadCmd_valid <= pkg_toStdLogic(false);
    if when_DataCache_l657 = '1' then
      dataReadCmd_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l657,io_cpu_execute_address)
  begin
    dataReadCmd_payload <= pkg_unsigned("XXXXXXXXX");
    if when_DataCache_l657 = '1' then
      dataReadCmd_payload <= pkg_extract(io_cpu_execute_address,10,2);
    end if;
  end process;

  process(when_DataCache_l843,when_DataCache_l1052,loader_done)
  begin
    tagsWriteCmd_valid <= pkg_toStdLogic(false);
    if when_DataCache_l843 = '1' then
      tagsWriteCmd_valid <= pkg_toStdLogic(true);
    end if;
    if when_DataCache_l1052 = '1' then
      tagsWriteCmd_valid <= pkg_toStdLogic(false);
    end if;
    if loader_done = '1' then
      tagsWriteCmd_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DataCache_l843,loader_done,loader_waysAllocator)
  begin
    tagsWriteCmd_payload_way <= pkg_stdLogicVector("XXXX");
    if when_DataCache_l843 = '1' then
      tagsWriteCmd_payload_way <= pkg_stdLogicVector("1111");
    end if;
    if loader_done = '1' then
      tagsWriteCmd_payload_way <= loader_waysAllocator;
    end if;
  end process;

  process(when_DataCache_l843,stageB_flusher_counter,loader_done,stageB_mmuRsp_physicalAddress)
  begin
    tagsWriteCmd_payload_address <= pkg_unsigned("XXXXXX");
    if when_DataCache_l843 = '1' then
      tagsWriteCmd_payload_address <= pkg_resize(stageB_flusher_counter,6);
    end if;
    if loader_done = '1' then
      tagsWriteCmd_payload_address <= pkg_extract(stageB_mmuRsp_physicalAddress,10,5);
    end if;
  end process;

  process(when_DataCache_l843,loader_done,loader_kill,loader_killReg)
  begin
    tagsWriteCmd_payload_data_valid <= 'X';
    if when_DataCache_l843 = '1' then
      tagsWriteCmd_payload_data_valid <= pkg_toStdLogic(false);
    end if;
    if loader_done = '1' then
      tagsWriteCmd_payload_data_valid <= (not (loader_kill or loader_killReg));
    end if;
  end process;

  process(loader_done,loader_error,io_mem_rsp_valid,io_mem_rsp_payload_error)
  begin
    tagsWriteCmd_payload_data_error <= 'X';
    if loader_done = '1' then
      tagsWriteCmd_payload_data_error <= (loader_error or (io_mem_rsp_valid and io_mem_rsp_payload_error));
    end if;
  end process;

  process(loader_done,stageB_mmuRsp_physicalAddress)
  begin
    tagsWriteCmd_payload_data_address <= pkg_unsigned("XXXXXXXXXXXXXXXXXXXXX");
    if loader_done = '1' then
      tagsWriteCmd_payload_data_address <= pkg_extract(stageB_mmuRsp_physicalAddress,31,11);
    end if;
  end process;

  process(stageB_cpuWriteToCache,when_DataCache_l912,when_DataCache_l1052,when_DataCache_l1076)
  begin
    dataWriteCmd_valid <= pkg_toStdLogic(false);
    if stageB_cpuWriteToCache = '1' then
      if when_DataCache_l912 = '1' then
        dataWriteCmd_valid <= pkg_toStdLogic(true);
      end if;
    end if;
    if when_DataCache_l1052 = '1' then
      dataWriteCmd_valid <= pkg_toStdLogic(false);
    end if;
    if when_DataCache_l1076 = '1' then
      dataWriteCmd_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(stageB_cpuWriteToCache,stageB_waysHits,when_DataCache_l1076,loader_waysAllocator)
  begin
    dataWriteCmd_payload_way <= pkg_stdLogicVector("XXXX");
    if stageB_cpuWriteToCache = '1' then
      dataWriteCmd_payload_way <= stageB_waysHits;
    end if;
    if when_DataCache_l1076 = '1' then
      dataWriteCmd_payload_way <= loader_waysAllocator;
    end if;
  end process;

  process(stageB_cpuWriteToCache,stageB_mmuRsp_physicalAddress,when_DataCache_l1076,loader_counter_value)
  begin
    dataWriteCmd_payload_address <= pkg_unsigned("XXXXXXXXX");
    if stageB_cpuWriteToCache = '1' then
      dataWriteCmd_payload_address <= pkg_extract(stageB_mmuRsp_physicalAddress,10,2);
    end if;
    if when_DataCache_l1076 = '1' then
      dataWriteCmd_payload_address <= unsigned(pkg_cat(std_logic_vector(pkg_extract(stageB_mmuRsp_physicalAddress,10,5)),std_logic_vector(loader_counter_value)));
    end if;
  end process;

  process(stageB_cpuWriteToCache,stageB_requestDataBypass,when_DataCache_l1076,io_mem_rsp_payload_data)
  begin
    dataWriteCmd_payload_data <= pkg_stdLogicVector("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
    if stageB_cpuWriteToCache = '1' then
      dataWriteCmd_payload_data(31 downto 0) <= stageB_requestDataBypass;
    end if;
    if when_DataCache_l1076 = '1' then
      dataWriteCmd_payload_data <= io_mem_rsp_payload_data;
    end if;
  end process;

  process(stageB_cpuWriteToCache,stageB_mask,when_DataCache_l1076)
  begin
    dataWriteCmd_payload_mask <= pkg_stdLogicVector("XXXX");
    if stageB_cpuWriteToCache = '1' then
      dataWriteCmd_payload_mask <= pkg_stdLogicVector("0000");
      if pkg_extract(pkg_unsigned("1"),0) = '1' then
        dataWriteCmd_payload_mask(3 downto 0) <= stageB_mask;
      end if;
    end if;
    if when_DataCache_l1076 = '1' then
      dataWriteCmd_payload_mask <= pkg_stdLogicVector("1111");
    end if;
  end process;

  when_DataCache_l657 <= (io_cpu_execute_isValid and (not io_cpu_memory_isStuck));
  process(when_DataCache_l843)
  begin
    io_cpu_execute_haltIt <= pkg_toStdLogic(false);
    if when_DataCache_l843 = '1' then
      io_cpu_execute_haltIt <= pkg_toStdLogic(true);
    end if;
  end process;

  rspSync <= pkg_toStdLogic(true);
  rspLast <= pkg_toStdLogic(true);
  io_mem_cmd_fire <= (io_mem_cmd_valid_read_buffer and io_mem_cmd_ready);
  when_DataCache_l679 <= (not io_cpu_writeBack_isStuck);
  process(io_cpu_execute_args_size)
  begin
    zz_stage0_mask <= pkg_stdLogicVector("XXXX");
    case io_cpu_execute_args_size is
      when "00" =>
        zz_stage0_mask <= pkg_stdLogicVector("0001");
      when "01" =>
        zz_stage0_mask <= pkg_stdLogicVector("0011");
      when "10" =>
        zz_stage0_mask <= pkg_stdLogicVector("1111");
      when others =>
    end case;
  end process;

  stage0_mask <= std_logic_vector(shift_left(unsigned(zz_stage0_mask),to_integer(pkg_extract(io_cpu_execute_address,1,0))));
  zz_stage0_dataColisions <= pkg_shiftRight(pkg_extract(io_cpu_execute_address,10,2),0);
  zz_stage0_dataColisions_1 <= pkg_extract(dataWriteCmd_payload_mask,3,0);
  process(dataWriteCmd_valid,dataWriteCmd_payload_way,dataWriteCmd_payload_address,zz_stage0_dataColisions,stage0_mask,zz_stage0_dataColisions_1)
  begin
    stage0_dataColisions(0) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,0)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stage0_dataColisions)) and pkg_toStdLogic((stage0_mask and zz_stage0_dataColisions_1) /= pkg_stdLogicVector("0000")));
    stage0_dataColisions(1) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,1)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stage0_dataColisions)) and pkg_toStdLogic((stage0_mask and zz_stage0_dataColisions_1) /= pkg_stdLogicVector("0000")));
    stage0_dataColisions(2) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,2)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stage0_dataColisions)) and pkg_toStdLogic((stage0_mask and zz_stage0_dataColisions_1) /= pkg_stdLogicVector("0000")));
    stage0_dataColisions(3) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,3)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stage0_dataColisions)) and pkg_toStdLogic((stage0_mask and zz_stage0_dataColisions_1) /= pkg_stdLogicVector("0000")));
  end process;

  stage0_wayInvalidate <= pkg_stdLogicVector("0000");
  stage0_isAmo <= pkg_toStdLogic(false);
  when_DataCache_l764 <= (not io_cpu_memory_isStuck);
  when_DataCache_l764_1 <= (not io_cpu_memory_isStuck);
  io_cpu_memory_isWrite <= stageA_request_wr;
  stageA_isAmo <= pkg_toStdLogic(false);
  stageA_isLrsc <= pkg_toStdLogic(false);
  stageA_wayHits <= pkg_cat(pkg_toStdLogicVector((pkg_toStdLogic(pkg_extract(io_cpu_memory_mmuRsp_physicalAddress,31,11) = ways_3_tagsReadRsp_address) and ways_3_tagsReadRsp_valid)),pkg_cat(pkg_toStdLogicVector((pkg_toStdLogic(pkg_extract(io_cpu_memory_mmuRsp_physicalAddress,31,11) = ways_2_tagsReadRsp_address) and ways_2_tagsReadRsp_valid)),pkg_cat(pkg_toStdLogicVector((pkg_toStdLogic(pkg_extract(io_cpu_memory_mmuRsp_physicalAddress,31,11) = ways_1_tagsReadRsp_address) and ways_1_tagsReadRsp_valid)),pkg_toStdLogicVector((pkg_toStdLogic(pkg_extract(io_cpu_memory_mmuRsp_physicalAddress,31,11) = ways_0_tagsReadRsp_address) and ways_0_tagsReadRsp_valid)))));
  when_DataCache_l764_2 <= (not io_cpu_memory_isStuck);
  when_DataCache_l764_3 <= (not io_cpu_memory_isStuck);
  zz_stageA_dataColisions_1 <= pkg_shiftRight(pkg_extract(io_cpu_memory_address,10,2),0);
  zz_stageA_dataColisions_2 <= pkg_extract(dataWriteCmd_payload_mask,3,0);
  process(dataWriteCmd_valid,dataWriteCmd_payload_way,dataWriteCmd_payload_address,zz_stageA_dataColisions_1,stageA_mask,zz_stageA_dataColisions_2)
  begin
    zz_stageA_dataColisions(0) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,0)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stageA_dataColisions_1)) and pkg_toStdLogic((stageA_mask and zz_stageA_dataColisions_2) /= pkg_stdLogicVector("0000")));
    zz_stageA_dataColisions(1) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,1)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stageA_dataColisions_1)) and pkg_toStdLogic((stageA_mask and zz_stageA_dataColisions_2) /= pkg_stdLogicVector("0000")));
    zz_stageA_dataColisions(2) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,2)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stageA_dataColisions_1)) and pkg_toStdLogic((stageA_mask and zz_stageA_dataColisions_2) /= pkg_stdLogicVector("0000")));
    zz_stageA_dataColisions(3) <= (((dataWriteCmd_valid and pkg_extract(dataWriteCmd_payload_way,3)) and pkg_toStdLogic(dataWriteCmd_payload_address = zz_stageA_dataColisions_1)) and pkg_toStdLogic((stageA_mask and zz_stageA_dataColisions_2) /= pkg_stdLogicVector("0000")));
  end process;

  stageA_dataColisions <= (stage0_dataColisions_regNextWhen or zz_stageA_dataColisions);
  when_DataCache_l815 <= (not io_cpu_writeBack_isStuck);
  process(when_DataCache_l1111)
  begin
    stageB_mmuRspFreeze <= pkg_toStdLogic(false);
    if when_DataCache_l1111 = '1' then
      stageB_mmuRspFreeze <= pkg_toStdLogic(true);
    end if;
  end process;

  when_DataCache_l817 <= ((not io_cpu_writeBack_isStuck) and (not stageB_mmuRspFreeze));
  when_DataCache_l814 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_1 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_2 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_3 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_4 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_5 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_6 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l814_7 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l813 <= (not io_cpu_writeBack_isStuck);
  stageB_consistancyHazard <= pkg_toStdLogic(false);
  when_DataCache_l813_1 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l813_2 <= (not io_cpu_writeBack_isStuck);
  when_DataCache_l813_3 <= (not io_cpu_writeBack_isStuck);
  stageB_waysHits <= (stageB_waysHitsBeforeInvalidate and pkg_not(stageB_wayInvalidate));
  stageB_waysHit <= pkg_toStdLogic(stageB_waysHits /= pkg_stdLogicVector("0000"));
  zz_stageB_dataMux <= pkg_extract(stageB_waysHits,3);
  zz_stageB_dataMux_1 <= (pkg_extract(stageB_waysHits,1) or zz_stageB_dataMux);
  zz_stageB_dataMux_2 <= (pkg_extract(stageB_waysHits,2) or zz_stageB_dataMux);
  stageB_dataMux <= zz_stageB_dataMux_3;
  when_DataCache_l813_4 <= (not io_cpu_writeBack_isStuck);
  process(io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l990,io_mem_cmd_ready,when_DataCache_l1052)
  begin
    stageB_loaderValid <= pkg_toStdLogic(false);
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '0' then
          if when_DataCache_l990 = '0' then
            if io_mem_cmd_ready = '1' then
              stageB_loaderValid <= pkg_toStdLogic(true);
            end if;
          end if;
        end if;
      end if;
    end if;
    if when_DataCache_l1052 = '1' then
      stageB_loaderValid <= pkg_toStdLogic(false);
    end if;
  end process;

  stageB_ioMemRspMuxed <= pkg_extract(io_mem_rsp_payload_data,31,0);
  process(io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l981,when_DataCache_l990,when_DataCache_l995,when_DataCache_l1052)
  begin
    io_cpu_writeBack_haltIt_read_buffer <= pkg_toStdLogic(true);
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '1' then
          if when_DataCache_l981 = '1' then
            io_cpu_writeBack_haltIt_read_buffer <= pkg_toStdLogic(false);
          end if;
        else
          if when_DataCache_l990 = '1' then
            if when_DataCache_l995 = '1' then
              io_cpu_writeBack_haltIt_read_buffer <= pkg_toStdLogic(false);
            end if;
          end if;
        end if;
      end if;
    end if;
    if when_DataCache_l1052 = '1' then
      io_cpu_writeBack_haltIt_read_buffer <= pkg_toStdLogic(false);
    end if;
  end process;

  stageB_flusher_hold <= pkg_toStdLogic(false);
  when_DataCache_l843 <= (not pkg_extract(stageB_flusher_counter,6));
  when_DataCache_l849 <= (not stageB_flusher_hold);
  io_cpu_flush_ready_read_buffer <= (stageB_flusher_waitDone and pkg_extract(stageB_flusher_counter,6));
  stageB_isAmo <= pkg_toStdLogic(false);
  stageB_isAmoCached <= pkg_toStdLogic(false);
  stageB_isExternalLsrc <= pkg_toStdLogic(false);
  stageB_isExternalAmo <= pkg_toStdLogic(false);
  stageB_requestDataBypass <= io_cpu_writeBack_storeData;
  process(io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l990)
  begin
    stageB_cpuWriteToCache <= pkg_toStdLogic(false);
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '0' then
          if when_DataCache_l990 = '1' then
            stageB_cpuWriteToCache <= pkg_toStdLogic(true);
          end if;
        end if;
      end if;
    end if;
  end process;

  when_DataCache_l912 <= (stageB_request_wr and stageB_waysHit);
  stageB_badPermissions <= (((not stageB_mmuRsp_allowWrite) and stageB_request_wr) or ((not stageB_mmuRsp_allowRead) and ((not stageB_request_wr) or stageB_isAmo)));
  stageB_loadStoreFault <= (io_cpu_writeBack_isValid and (stageB_mmuRsp_exception or stageB_badPermissions));
  process(io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l990,when_DataCache_l1006,when_DataCache_l1061,when_DataCache_l1108)
  begin
    io_cpu_redo_read_buffer <= pkg_toStdLogic(false);
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '0' then
          if when_DataCache_l990 = '1' then
            if when_DataCache_l1006 = '1' then
              io_cpu_redo_read_buffer <= pkg_toStdLogic(true);
            end if;
          end if;
        end if;
      end if;
    end if;
    if when_DataCache_l1061 = '1' then
      io_cpu_redo_read_buffer <= pkg_toStdLogic(true);
    end if;
    if when_DataCache_l1108 = '1' then
      io_cpu_redo_read_buffer <= pkg_toStdLogic(true);
    end if;
  end process;

  process(stageB_bypassCache,stageB_request_wr,io_mem_rsp_valid,io_mem_rsp_payload_error,stageB_waysHits,stageB_tagsReadRsp_3_error,stageB_tagsReadRsp_2_error,stageB_tagsReadRsp_1_error,stageB_tagsReadRsp_0_error,stageB_loadStoreFault,stageB_mmuRsp_isPaging)
  begin
    io_cpu_writeBack_accessError_read_buffer <= pkg_toStdLogic(false);
    if stageB_bypassCache = '1' then
      io_cpu_writeBack_accessError_read_buffer <= ((((not stageB_request_wr) and pkg_toStdLogic(true)) and io_mem_rsp_valid) and io_mem_rsp_payload_error);
    else
      io_cpu_writeBack_accessError_read_buffer <= (pkg_toStdLogic((stageB_waysHits and pkg_cat(pkg_toStdLogicVector(stageB_tagsReadRsp_3_error),pkg_cat(pkg_toStdLogicVector(stageB_tagsReadRsp_2_error),pkg_cat(pkg_toStdLogicVector(stageB_tagsReadRsp_1_error),pkg_toStdLogicVector(stageB_tagsReadRsp_0_error))))) /= pkg_stdLogicVector("0000")) or (stageB_loadStoreFault and (not stageB_mmuRsp_isPaging)));
    end if;
  end process;

  io_cpu_writeBack_mmuException_read_buffer <= (stageB_loadStoreFault and stageB_mmuRsp_isPaging);
  io_cpu_writeBack_unalignedAccess_read_buffer <= (io_cpu_writeBack_isValid and stageB_unaligned);
  io_cpu_writeBack_isWrite <= stageB_request_wr;
  process(io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,memCmdSent,when_DataCache_l990,stageB_request_wr,when_DataCache_l1018,when_DataCache_l1052)
  begin
    io_mem_cmd_valid_read_buffer <= pkg_toStdLogic(false);
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '1' then
          io_mem_cmd_valid_read_buffer <= (not memCmdSent);
        else
          if when_DataCache_l990 = '1' then
            if stageB_request_wr = '1' then
              io_mem_cmd_valid_read_buffer <= pkg_toStdLogic(true);
            end if;
          else
            if when_DataCache_l1018 = '1' then
              io_mem_cmd_valid_read_buffer <= pkg_toStdLogic(true);
            end if;
          end if;
        end if;
      end if;
    end if;
    if when_DataCache_l1052 = '1' then
      io_mem_cmd_valid_read_buffer <= pkg_toStdLogic(false);
    end if;
  end process;

  process(stageB_mmuRsp_physicalAddress,io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l990)
  begin
    io_mem_cmd_payload_address <= stageB_mmuRsp_physicalAddress;
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '0' then
          if when_DataCache_l990 = '0' then
            io_mem_cmd_payload_address(4 downto 0) <= pkg_unsigned("00000");
          end if;
        end if;
      end if;
    end if;
  end process;

  io_mem_cmd_payload_last <= pkg_toStdLogic(true);
  process(stageB_request_wr,io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l990)
  begin
    io_mem_cmd_payload_wr <= stageB_request_wr;
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '0' then
          if when_DataCache_l990 = '0' then
            io_mem_cmd_payload_wr <= pkg_toStdLogic(false);
          end if;
        end if;
      end if;
    end if;
  end process;

  io_mem_cmd_payload_mask <= stageB_mask;
  io_mem_cmd_payload_data <= stageB_requestDataBypass;
  io_mem_cmd_payload_uncached <= stageB_mmuRsp_isIoAccess;
  process(stageB_request_size,io_cpu_writeBack_isValid,stageB_isExternalAmo,when_DataCache_l977,when_DataCache_l990)
  begin
    io_mem_cmd_payload_size <= pkg_resize(stageB_request_size,3);
    if io_cpu_writeBack_isValid = '1' then
      if stageB_isExternalAmo = '0' then
        if when_DataCache_l977 = '0' then
          if when_DataCache_l990 = '0' then
            io_mem_cmd_payload_size <= pkg_unsigned("101");
          end if;
        end if;
      end if;
    end if;
  end process;

  stageB_bypassCache <= ((stageB_mmuRsp_isIoAccess or stageB_isExternalLsrc) or stageB_isExternalAmo);
  io_cpu_writeBack_keepMemRspData <= pkg_toStdLogic(false);
  when_DataCache_l981 <= pkg_mux((not stageB_request_wr),(io_mem_rsp_valid and rspSync),io_mem_cmd_ready);
  when_DataCache_l990 <= (stageB_waysHit or (stageB_request_wr and (not stageB_isAmoCached)));
  when_DataCache_l995 <= ((not stageB_request_wr) or io_mem_cmd_ready);
  when_DataCache_l1006 <= (((not stageB_request_wr) or stageB_isAmoCached) and pkg_toStdLogic((stageB_dataColisions and stageB_waysHits) /= pkg_stdLogicVector("0000")));
  when_DataCache_l1018 <= (not memCmdSent);
  when_DataCache_l977 <= (stageB_mmuRsp_isIoAccess or stageB_isExternalLsrc);
  process(stageB_bypassCache,stageB_ioMemRspMuxed,stageB_dataMux)
  begin
    if stageB_bypassCache = '1' then
      io_cpu_writeBack_data <= stageB_ioMemRspMuxed;
    else
      io_cpu_writeBack_data <= stageB_dataMux;
    end if;
  end process;

  when_DataCache_l1052 <= ((((stageB_consistancyHazard or stageB_mmuRsp_refilling) or io_cpu_writeBack_accessError_read_buffer) or io_cpu_writeBack_mmuException_read_buffer) or io_cpu_writeBack_unalignedAccess_read_buffer);
  when_DataCache_l1061 <= (io_cpu_writeBack_isValid and (stageB_mmuRsp_refilling or stageB_consistancyHazard));
  process(when_DataCache_l1076)
  begin
    loader_counter_willIncrement <= pkg_toStdLogic(false);
    if when_DataCache_l1076 = '1' then
      loader_counter_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  loader_counter_willClear <= pkg_toStdLogic(false);
  loader_counter_willOverflowIfInc <= pkg_toStdLogic(loader_counter_value = pkg_unsigned("111"));
  loader_counter_willOverflow <= (loader_counter_willOverflowIfInc and loader_counter_willIncrement);
  process(loader_counter_value,loader_counter_willIncrement,loader_counter_willClear)
  begin
    loader_counter_valueNext <= (loader_counter_value + pkg_resize(unsigned(pkg_toStdLogicVector(loader_counter_willIncrement)),3));
    if loader_counter_willClear = '1' then
      loader_counter_valueNext <= pkg_unsigned("000");
    end if;
  end process;

  loader_kill <= pkg_toStdLogic(false);
  when_DataCache_l1076 <= ((loader_valid and io_mem_rsp_valid) and rspLast);
  loader_done <= loader_counter_willOverflow;
  when_DataCache_l1104 <= (not loader_valid);
  when_DataCache_l1108 <= (loader_valid and (not loader_valid_regNext));
  io_cpu_execute_refilling <= loader_valid;
  when_DataCache_l1111 <= (stageB_loaderValid or loader_valid);
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      tagsWriteLastCmd_valid <= tagsWriteCmd_valid;
      tagsWriteLastCmd_payload_way <= tagsWriteCmd_payload_way;
      tagsWriteLastCmd_payload_address <= tagsWriteCmd_payload_address;
      tagsWriteLastCmd_payload_data_valid <= tagsWriteCmd_payload_data_valid;
      tagsWriteLastCmd_payload_data_error <= tagsWriteCmd_payload_data_error;
      tagsWriteLastCmd_payload_data_address <= tagsWriteCmd_payload_data_address;
      if when_DataCache_l764 = '1' then
        stageA_request_wr <= io_cpu_execute_args_wr;
        stageA_request_size <= io_cpu_execute_args_size;
        stageA_request_totalyConsistent <= io_cpu_execute_args_totalyConsistent;
      end if;
      if when_DataCache_l764_1 = '1' then
        stageA_mask <= stage0_mask;
      end if;
      if when_DataCache_l764_2 = '1' then
        stageA_wayInvalidate <= stage0_wayInvalidate;
      end if;
      if when_DataCache_l764_3 = '1' then
        stage0_dataColisions_regNextWhen <= stage0_dataColisions;
      end if;
      if when_DataCache_l815 = '1' then
        stageB_request_wr <= stageA_request_wr;
        stageB_request_size <= stageA_request_size;
        stageB_request_totalyConsistent <= stageA_request_totalyConsistent;
      end if;
      if when_DataCache_l817 = '1' then
        stageB_mmuRsp_physicalAddress <= io_cpu_memory_mmuRsp_physicalAddress;
        stageB_mmuRsp_isIoAccess <= io_cpu_memory_mmuRsp_isIoAccess;
        stageB_mmuRsp_isPaging <= io_cpu_memory_mmuRsp_isPaging;
        stageB_mmuRsp_allowRead <= io_cpu_memory_mmuRsp_allowRead;
        stageB_mmuRsp_allowWrite <= io_cpu_memory_mmuRsp_allowWrite;
        stageB_mmuRsp_allowExecute <= io_cpu_memory_mmuRsp_allowExecute;
        stageB_mmuRsp_exception <= io_cpu_memory_mmuRsp_exception;
        stageB_mmuRsp_refilling <= io_cpu_memory_mmuRsp_refilling;
        stageB_mmuRsp_bypassTranslation <= io_cpu_memory_mmuRsp_bypassTranslation;
      end if;
      if when_DataCache_l814 = '1' then
        stageB_tagsReadRsp_0_valid <= ways_0_tagsReadRsp_valid;
        stageB_tagsReadRsp_0_error <= ways_0_tagsReadRsp_error;
        stageB_tagsReadRsp_0_address <= ways_0_tagsReadRsp_address;
      end if;
      if when_DataCache_l814_1 = '1' then
        stageB_tagsReadRsp_1_valid <= ways_1_tagsReadRsp_valid;
        stageB_tagsReadRsp_1_error <= ways_1_tagsReadRsp_error;
        stageB_tagsReadRsp_1_address <= ways_1_tagsReadRsp_address;
      end if;
      if when_DataCache_l814_2 = '1' then
        stageB_tagsReadRsp_2_valid <= ways_2_tagsReadRsp_valid;
        stageB_tagsReadRsp_2_error <= ways_2_tagsReadRsp_error;
        stageB_tagsReadRsp_2_address <= ways_2_tagsReadRsp_address;
      end if;
      if when_DataCache_l814_3 = '1' then
        stageB_tagsReadRsp_3_valid <= ways_3_tagsReadRsp_valid;
        stageB_tagsReadRsp_3_error <= ways_3_tagsReadRsp_error;
        stageB_tagsReadRsp_3_address <= ways_3_tagsReadRsp_address;
      end if;
      if when_DataCache_l814_4 = '1' then
        stageB_dataReadRsp_0 <= ways_0_dataReadRsp;
      end if;
      if when_DataCache_l814_5 = '1' then
        stageB_dataReadRsp_1 <= ways_1_dataReadRsp;
      end if;
      if when_DataCache_l814_6 = '1' then
        stageB_dataReadRsp_2 <= ways_2_dataReadRsp;
      end if;
      if when_DataCache_l814_7 = '1' then
        stageB_dataReadRsp_3 <= ways_3_dataReadRsp;
      end if;
      if when_DataCache_l813 = '1' then
        stageB_wayInvalidate <= stageA_wayInvalidate;
      end if;
      if when_DataCache_l813_1 = '1' then
        stageB_dataColisions <= stageA_dataColisions;
      end if;
      if when_DataCache_l813_2 = '1' then
        stageB_unaligned <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector((pkg_toStdLogic(stageA_request_size = pkg_unsigned("10")) and pkg_toStdLogic(pkg_extract(io_cpu_memory_address,1,0) /= pkg_unsigned("00")))),pkg_toStdLogicVector((pkg_toStdLogic(stageA_request_size = pkg_unsigned("01")) and pkg_toStdLogic(pkg_extract(io_cpu_memory_address,0,0) /= pkg_unsigned("0"))))) /= pkg_stdLogicVector("00"));
      end if;
      if when_DataCache_l813_3 = '1' then
        stageB_waysHitsBeforeInvalidate <= stageA_wayHits;
      end if;
      if when_DataCache_l813_4 = '1' then
        stageB_mask <= stageA_mask;
      end if;
      loader_valid_regNext <= loader_valid;
    end if;
  end process;

  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      memCmdSent <= pkg_toStdLogic(false);
      stageB_flusher_waitDone <= pkg_toStdLogic(false);
      stageB_flusher_counter <= pkg_unsigned("0000000");
      stageB_flusher_start <= pkg_toStdLogic(true);
      loader_valid <= pkg_toStdLogic(false);
      loader_counter_value <= pkg_unsigned("000");
      loader_waysAllocator <= pkg_stdLogicVector("0001");
      loader_error <= pkg_toStdLogic(false);
      loader_killReg <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if io_mem_cmd_fire = '1' then
        memCmdSent <= pkg_toStdLogic(true);
      end if;
      if when_DataCache_l679 = '1' then
        memCmdSent <= pkg_toStdLogic(false);
      end if;
      if io_cpu_flush_ready_read_buffer = '1' then
        stageB_flusher_waitDone <= pkg_toStdLogic(false);
      end if;
      if when_DataCache_l843 = '1' then
        if when_DataCache_l849 = '1' then
          stageB_flusher_counter <= (stageB_flusher_counter + pkg_unsigned("0000001"));
        end if;
      end if;
      stageB_flusher_start <= (((((((not stageB_flusher_waitDone) and (not stageB_flusher_start)) and io_cpu_flush_valid) and (not io_cpu_execute_isValid)) and (not io_cpu_memory_isValid)) and (not io_cpu_writeBack_isValid)) and (not io_cpu_redo_read_buffer));
      if stageB_flusher_start = '1' then
        stageB_flusher_waitDone <= pkg_toStdLogic(true);
        stageB_flusher_counter <= pkg_unsigned("0000000");
      end if;
      assert (not ((io_cpu_writeBack_isValid and (not io_cpu_writeBack_haltIt_read_buffer)) and io_cpu_writeBack_isStuck)) = '1' report "writeBack stuck by another plugin is not allowed"  severity ERROR;
      if stageB_loaderValid = '1' then
        loader_valid <= pkg_toStdLogic(true);
      end if;
      loader_counter_value <= loader_counter_valueNext;
      if loader_kill = '1' then
        loader_killReg <= pkg_toStdLogic(true);
      end if;
      if when_DataCache_l1076 = '1' then
        loader_error <= (loader_error or io_mem_rsp_payload_error);
      end if;
      if loader_done = '1' then
        loader_valid <= pkg_toStdLogic(false);
        loader_error <= pkg_toStdLogic(false);
        loader_killReg <= pkg_toStdLogic(false);
      end if;
      if when_DataCache_l1104 = '1' then
        loader_waysAllocator <= pkg_resize(pkg_cat(loader_waysAllocator,pkg_toStdLogicVector(pkg_extract(loader_waysAllocator,3))),4);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity FlowCCByToggle is
  port(
    io_input_valid : in std_logic;
    io_input_payload_last : in std_logic;
    io_input_payload_fragment : in std_logic_vector(0 downto 0);
    io_output_valid : out std_logic;
    io_output_payload_last : out std_logic;
    io_output_payload_fragment : out std_logic_vector(0 downto 0);
    TCK : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_systemReset : in std_logic
  );
end FlowCCByToggle;

architecture arch of FlowCCByToggle is
  signal inputArea_target_buffercc_io_dataOut : std_logic;

  signal outHitSignal : std_logic;
  signal inputArea_target : std_logic := '0';
  signal inputArea_data_last : std_logic;
  signal inputArea_data_fragment : std_logic_vector(0 downto 0);
  signal outputArea_target : std_logic;
  signal outputArea_hit : std_logic;
  signal outputArea_flow_valid : std_logic;
  signal outputArea_flow_payload_last : std_logic;
  signal outputArea_flow_payload_fragment : std_logic_vector(0 downto 0);
  signal outputArea_flow_m2sPipe_valid : std_logic;
  signal outputArea_flow_m2sPipe_payload_last : std_logic;
  signal outputArea_flow_m2sPipe_payload_fragment : std_logic_vector(0 downto 0);
begin
  inputArea_target_buffercc : entity work.BufferCC_1
    port map ( 
      io_dataIn => inputArea_target,
      io_dataOut => inputArea_target_buffercc_io_dataOut,
      io_mainClk => io_mainClk,
      resetCtrl_systemReset => resetCtrl_systemReset 
    );
  outputArea_target <= inputArea_target_buffercc_io_dataOut;
  outputArea_flow_valid <= pkg_toStdLogic(outputArea_target /= outputArea_hit);
  outputArea_flow_payload_last <= inputArea_data_last;
  outputArea_flow_payload_fragment <= inputArea_data_fragment;
  io_output_valid <= outputArea_flow_m2sPipe_valid;
  io_output_payload_last <= outputArea_flow_m2sPipe_payload_last;
  io_output_payload_fragment <= outputArea_flow_m2sPipe_payload_fragment;
  process(TCK)
  begin
    if rising_edge(TCK) then
      if io_input_valid = '1' then
        inputArea_target <= (not inputArea_target);
        inputArea_data_last <= io_input_payload_last;
        inputArea_data_fragment <= io_input_payload_fragment;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      outputArea_hit <= outputArea_target;
      if outputArea_flow_valid = '1' then
        outputArea_flow_m2sPipe_payload_last <= outputArea_flow_payload_last;
        outputArea_flow_m2sPipe_payload_fragment <= outputArea_flow_payload_fragment;
      end if;
    end if;
  end process;

  process(io_mainClk, resetCtrl_systemReset)
  begin
    if resetCtrl_systemReset = '1' then
      outputArea_flow_m2sPipe_valid <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      outputArea_flow_m2sPipe_valid <= outputArea_flow_valid;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4ReadOnlyErrorSlave is
  port(
    io_axi_ar_valid : in std_logic;
    io_axi_ar_ready : out std_logic;
    io_axi_ar_payload_addr : in unsigned(31 downto 0);
    io_axi_ar_payload_len : in unsigned(7 downto 0);
    io_axi_ar_payload_burst : in std_logic_vector(1 downto 0);
    io_axi_ar_payload_cache : in std_logic_vector(3 downto 0);
    io_axi_ar_payload_prot : in std_logic_vector(2 downto 0);
    io_axi_r_valid : out std_logic;
    io_axi_r_ready : in std_logic;
    io_axi_r_payload_data : out std_logic_vector(31 downto 0);
    io_axi_r_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_payload_last : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4ReadOnlyErrorSlave;

architecture arch of Axi4ReadOnlyErrorSlave is
  signal io_axi_ar_ready_read_buffer : std_logic;

  signal sendRsp : std_logic;
  signal remaining : unsigned(7 downto 0);
  signal remainingZero : std_logic;
  signal io_axi_ar_fire : std_logic;
begin
  io_axi_ar_ready <= io_axi_ar_ready_read_buffer;
  remainingZero <= pkg_toStdLogic(remaining = pkg_unsigned("00000000"));
  io_axi_ar_ready_read_buffer <= (not sendRsp);
  io_axi_ar_fire <= (io_axi_ar_valid and io_axi_ar_ready_read_buffer);
  io_axi_r_valid <= sendRsp;
  io_axi_r_payload_resp <= pkg_stdLogicVector("11");
  io_axi_r_payload_last <= remainingZero;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      sendRsp <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if io_axi_ar_fire = '1' then
        sendRsp <= pkg_toStdLogic(true);
      end if;
      if sendRsp = '1' then
        if io_axi_r_ready = '1' then
          if remainingZero = '1' then
            sendRsp <= pkg_toStdLogic(false);
          end if;
        end if;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_axi_ar_fire = '1' then
        remaining <= io_axi_ar_payload_len;
      end if;
      if sendRsp = '1' then
        if io_axi_r_ready = '1' then
          remaining <= (remaining - pkg_unsigned("00000001"));
        end if;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4SharedErrorSlave is
  port(
    io_axi_arw_valid : in std_logic;
    io_axi_arw_ready : out std_logic;
    io_axi_arw_payload_addr : in unsigned(31 downto 0);
    io_axi_arw_payload_len : in unsigned(7 downto 0);
    io_axi_arw_payload_size : in unsigned(2 downto 0);
    io_axi_arw_payload_cache : in std_logic_vector(3 downto 0);
    io_axi_arw_payload_prot : in std_logic_vector(2 downto 0);
    io_axi_arw_payload_write : in std_logic;
    io_axi_w_valid : in std_logic;
    io_axi_w_ready : out std_logic;
    io_axi_w_payload_data : in std_logic_vector(31 downto 0);
    io_axi_w_payload_strb : in std_logic_vector(3 downto 0);
    io_axi_w_payload_last : in std_logic;
    io_axi_b_valid : out std_logic;
    io_axi_b_ready : in std_logic;
    io_axi_b_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_valid : out std_logic;
    io_axi_r_ready : in std_logic;
    io_axi_r_payload_data : out std_logic_vector(31 downto 0);
    io_axi_r_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_payload_last : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4SharedErrorSlave;

architecture arch of Axi4SharedErrorSlave is
  signal io_axi_arw_ready_read_buffer : std_logic;
  signal io_axi_w_ready_read_buffer : std_logic;
  signal io_axi_b_valid_read_buffer : std_logic;

  signal consumeData : std_logic;
  signal sendReadRsp : std_logic;
  signal sendWriteRsp : std_logic;
  signal remaining : unsigned(7 downto 0);
  signal remainingZero : std_logic;
  signal io_axi_arw_fire : std_logic;
  signal io_axi_w_fire : std_logic;
  signal when_Axi4ErrorSlave_l92 : std_logic;
  signal io_axi_b_fire : std_logic;
begin
  io_axi_arw_ready <= io_axi_arw_ready_read_buffer;
  io_axi_w_ready <= io_axi_w_ready_read_buffer;
  io_axi_b_valid <= io_axi_b_valid_read_buffer;
  remainingZero <= pkg_toStdLogic(remaining = pkg_unsigned("00000000"));
  io_axi_arw_ready_read_buffer <= (not ((consumeData or sendWriteRsp) or sendReadRsp));
  io_axi_arw_fire <= (io_axi_arw_valid and io_axi_arw_ready_read_buffer);
  io_axi_w_ready_read_buffer <= consumeData;
  io_axi_w_fire <= (io_axi_w_valid and io_axi_w_ready_read_buffer);
  when_Axi4ErrorSlave_l92 <= (io_axi_w_fire and io_axi_w_payload_last);
  io_axi_b_valid_read_buffer <= sendWriteRsp;
  io_axi_b_payload_resp <= pkg_stdLogicVector("11");
  io_axi_b_fire <= (io_axi_b_valid_read_buffer and io_axi_b_ready);
  io_axi_r_valid <= sendReadRsp;
  io_axi_r_payload_resp <= pkg_stdLogicVector("11");
  io_axi_r_payload_last <= remainingZero;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      consumeData <= pkg_toStdLogic(false);
      sendReadRsp <= pkg_toStdLogic(false);
      sendWriteRsp <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if io_axi_arw_fire = '1' then
        consumeData <= io_axi_arw_payload_write;
        sendReadRsp <= (not io_axi_arw_payload_write);
      end if;
      if when_Axi4ErrorSlave_l92 = '1' then
        consumeData <= pkg_toStdLogic(false);
        sendWriteRsp <= pkg_toStdLogic(true);
      end if;
      if io_axi_b_fire = '1' then
        sendWriteRsp <= pkg_toStdLogic(false);
      end if;
      if sendReadRsp = '1' then
        if io_axi_r_ready = '1' then
          if remainingZero = '1' then
            sendReadRsp <= pkg_toStdLogic(false);
          end if;
        end if;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_axi_arw_fire = '1' then
        remaining <= io_axi_arw_payload_len;
      end if;
      if sendReadRsp = '1' then
        if io_axi_r_ready = '1' then
          remaining <= (remaining - pkg_unsigned("00000001"));
        end if;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamArbiter is
  port(
    io_inputs_0_valid : in std_logic;
    io_inputs_0_ready : out std_logic;
    io_inputs_0_payload_addr : in unsigned(14 downto 0);
    io_inputs_0_payload_id : in unsigned(2 downto 0);
    io_inputs_0_payload_len : in unsigned(7 downto 0);
    io_inputs_0_payload_size : in unsigned(2 downto 0);
    io_inputs_0_payload_burst : in std_logic_vector(1 downto 0);
    io_inputs_0_payload_write : in std_logic;
    io_inputs_1_valid : in std_logic;
    io_inputs_1_ready : out std_logic;
    io_inputs_1_payload_addr : in unsigned(14 downto 0);
    io_inputs_1_payload_id : in unsigned(2 downto 0);
    io_inputs_1_payload_len : in unsigned(7 downto 0);
    io_inputs_1_payload_size : in unsigned(2 downto 0);
    io_inputs_1_payload_burst : in std_logic_vector(1 downto 0);
    io_inputs_1_payload_write : in std_logic;
    io_output_valid : out std_logic;
    io_output_ready : in std_logic;
    io_output_payload_addr : out unsigned(14 downto 0);
    io_output_payload_id : out unsigned(2 downto 0);
    io_output_payload_len : out unsigned(7 downto 0);
    io_output_payload_size : out unsigned(2 downto 0);
    io_output_payload_burst : out std_logic_vector(1 downto 0);
    io_output_payload_write : out std_logic;
    io_chosen : out unsigned(0 downto 0);
    io_chosenOH : out std_logic_vector(1 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamArbiter;

architecture arch of StreamArbiter is
  signal io_output_valid_read_buffer : std_logic;
  signal io_chosenOH_read_buffer : std_logic_vector(1 downto 0);

  signal locked : std_logic;
  signal maskProposal_0 : std_logic;
  signal maskProposal_1 : std_logic;
  signal maskLocked_0 : std_logic;
  signal maskLocked_1 : std_logic;
  signal maskRouted_0 : std_logic;
  signal maskRouted_1 : std_logic;
  signal zz_maskProposal_0 : unsigned(1 downto 0);
  signal zz_maskProposal_0_1 : unsigned(3 downto 0);
  signal zz_maskProposal_0_2 : unsigned(3 downto 0);
  signal zz_maskProposal_0_3 : std_logic_vector(1 downto 0);
  signal io_output_fire : std_logic;
  signal zz_io_chosen : std_logic;
begin
  io_output_valid <= io_output_valid_read_buffer;
  io_chosenOH <= io_chosenOH_read_buffer;
  maskRouted_0 <= pkg_mux(locked,maskLocked_0,maskProposal_0);
  maskRouted_1 <= pkg_mux(locked,maskLocked_1,maskProposal_1);
  zz_maskProposal_0 <= unsigned(pkg_cat(pkg_toStdLogicVector(io_inputs_1_valid),pkg_toStdLogicVector(io_inputs_0_valid)));
  zz_maskProposal_0_1 <= unsigned(pkg_cat(std_logic_vector(zz_maskProposal_0),std_logic_vector(zz_maskProposal_0)));
  zz_maskProposal_0_2 <= (zz_maskProposal_0_1 and pkg_not((zz_maskProposal_0_1 - pkg_resize(unsigned(pkg_cat(pkg_toStdLogicVector(maskLocked_0),pkg_toStdLogicVector(maskLocked_1))),4))));
  zz_maskProposal_0_3 <= std_logic_vector((pkg_extract(zz_maskProposal_0_2,3,2) or pkg_extract(zz_maskProposal_0_2,1,0)));
  maskProposal_0 <= pkg_extract(zz_maskProposal_0_3,0);
  maskProposal_1 <= pkg_extract(zz_maskProposal_0_3,1);
  io_output_fire <= (io_output_valid_read_buffer and io_output_ready);
  io_output_valid_read_buffer <= ((io_inputs_0_valid and maskRouted_0) or (io_inputs_1_valid and maskRouted_1));
  io_output_payload_addr <= pkg_mux(maskRouted_0,io_inputs_0_payload_addr,io_inputs_1_payload_addr);
  io_output_payload_id <= pkg_mux(maskRouted_0,io_inputs_0_payload_id,io_inputs_1_payload_id);
  io_output_payload_len <= pkg_mux(maskRouted_0,io_inputs_0_payload_len,io_inputs_1_payload_len);
  io_output_payload_size <= pkg_mux(maskRouted_0,io_inputs_0_payload_size,io_inputs_1_payload_size);
  io_output_payload_burst <= pkg_mux(maskRouted_0,io_inputs_0_payload_burst,io_inputs_1_payload_burst);
  io_output_payload_write <= pkg_mux(maskRouted_0,io_inputs_0_payload_write,io_inputs_1_payload_write);
  io_inputs_0_ready <= (maskRouted_0 and io_output_ready);
  io_inputs_1_ready <= (maskRouted_1 and io_output_ready);
  io_chosenOH_read_buffer <= pkg_cat(pkg_toStdLogicVector(maskRouted_1),pkg_toStdLogicVector(maskRouted_0));
  zz_io_chosen <= pkg_extract(io_chosenOH_read_buffer,1);
  io_chosen <= unsigned(pkg_toStdLogicVector(zz_io_chosen));
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      locked <= pkg_toStdLogic(false);
      maskLocked_0 <= pkg_toStdLogic(false);
      maskLocked_1 <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      if io_output_valid_read_buffer = '1' then
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end if;
      if io_output_valid_read_buffer = '1' then
        locked <= pkg_toStdLogic(true);
      end if;
      if io_output_fire = '1' then
        locked <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamFork is
  port(
    io_input_valid : in std_logic;
    io_input_ready : out std_logic;
    io_input_payload_addr : in unsigned(14 downto 0);
    io_input_payload_id : in unsigned(2 downto 0);
    io_input_payload_len : in unsigned(7 downto 0);
    io_input_payload_size : in unsigned(2 downto 0);
    io_input_payload_burst : in std_logic_vector(1 downto 0);
    io_input_payload_write : in std_logic;
    io_outputs_0_valid : out std_logic;
    io_outputs_0_ready : in std_logic;
    io_outputs_0_payload_addr : out unsigned(14 downto 0);
    io_outputs_0_payload_id : out unsigned(2 downto 0);
    io_outputs_0_payload_len : out unsigned(7 downto 0);
    io_outputs_0_payload_size : out unsigned(2 downto 0);
    io_outputs_0_payload_burst : out std_logic_vector(1 downto 0);
    io_outputs_0_payload_write : out std_logic;
    io_outputs_1_valid : out std_logic;
    io_outputs_1_ready : in std_logic;
    io_outputs_1_payload_addr : out unsigned(14 downto 0);
    io_outputs_1_payload_id : out unsigned(2 downto 0);
    io_outputs_1_payload_len : out unsigned(7 downto 0);
    io_outputs_1_payload_size : out unsigned(2 downto 0);
    io_outputs_1_payload_burst : out std_logic_vector(1 downto 0);
    io_outputs_1_payload_write : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamFork;

architecture arch of StreamFork is
  signal io_outputs_0_valid_read_buffer : std_logic;
  signal io_outputs_1_valid_read_buffer : std_logic;
  signal io_input_ready_read_buffer : std_logic;

  signal zz_io_outputs_0_valid : std_logic;
  signal zz_io_outputs_1_valid : std_logic;
  signal when_Stream_l817 : std_logic;
  signal when_Stream_l817_1 : std_logic;
  signal io_outputs_0_fire : std_logic;
  signal io_outputs_1_fire : std_logic;
begin
  io_outputs_0_valid <= io_outputs_0_valid_read_buffer;
  io_outputs_1_valid <= io_outputs_1_valid_read_buffer;
  io_input_ready <= io_input_ready_read_buffer;
  process(when_Stream_l817,when_Stream_l817_1)
  begin
    io_input_ready_read_buffer <= pkg_toStdLogic(true);
    if when_Stream_l817 = '1' then
      io_input_ready_read_buffer <= pkg_toStdLogic(false);
    end if;
    if when_Stream_l817_1 = '1' then
      io_input_ready_read_buffer <= pkg_toStdLogic(false);
    end if;
  end process;

  when_Stream_l817 <= ((not io_outputs_0_ready) and zz_io_outputs_0_valid);
  when_Stream_l817_1 <= ((not io_outputs_1_ready) and zz_io_outputs_1_valid);
  io_outputs_0_valid_read_buffer <= (io_input_valid and zz_io_outputs_0_valid);
  io_outputs_0_payload_addr <= io_input_payload_addr;
  io_outputs_0_payload_id <= io_input_payload_id;
  io_outputs_0_payload_len <= io_input_payload_len;
  io_outputs_0_payload_size <= io_input_payload_size;
  io_outputs_0_payload_burst <= io_input_payload_burst;
  io_outputs_0_payload_write <= io_input_payload_write;
  io_outputs_0_fire <= (io_outputs_0_valid_read_buffer and io_outputs_0_ready);
  io_outputs_1_valid_read_buffer <= (io_input_valid and zz_io_outputs_1_valid);
  io_outputs_1_payload_addr <= io_input_payload_addr;
  io_outputs_1_payload_id <= io_input_payload_id;
  io_outputs_1_payload_len <= io_input_payload_len;
  io_outputs_1_payload_size <= io_input_payload_size;
  io_outputs_1_payload_burst <= io_input_payload_burst;
  io_outputs_1_payload_write <= io_input_payload_write;
  io_outputs_1_fire <= (io_outputs_1_valid_read_buffer and io_outputs_1_ready);
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      zz_io_outputs_0_valid <= pkg_toStdLogic(true);
      zz_io_outputs_1_valid <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      if io_outputs_0_fire = '1' then
        zz_io_outputs_0_valid <= pkg_toStdLogic(false);
      end if;
      if io_outputs_1_fire = '1' then
        zz_io_outputs_1_valid <= pkg_toStdLogic(false);
      end if;
      if io_input_ready_read_buffer = '1' then
        zz_io_outputs_0_valid <= pkg_toStdLogic(true);
        zz_io_outputs_1_valid <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamFifoLowLatency is
  port(
    io_push_valid : in std_logic;
    io_push_ready : out std_logic;
    io_pop_valid : out std_logic;
    io_pop_ready : in std_logic;
    io_flush : in std_logic;
    io_occupancy : out unsigned(2 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamFifoLowLatency;

architecture arch of StreamFifoLowLatency is
  signal io_push_ready_read_buffer : std_logic;
  signal io_pop_valid_read_buffer : std_logic;

  signal pushPtr_willIncrement : std_logic;
  signal pushPtr_willClear : std_logic;
  signal pushPtr_valueNext : unsigned(1 downto 0);
  signal pushPtr_value : unsigned(1 downto 0);
  signal pushPtr_willOverflowIfInc : std_logic;
  signal pushPtr_willOverflow : std_logic;
  signal popPtr_willIncrement : std_logic;
  signal popPtr_willClear : std_logic;
  signal popPtr_valueNext : unsigned(1 downto 0);
  signal popPtr_value : unsigned(1 downto 0);
  signal popPtr_willOverflowIfInc : std_logic;
  signal popPtr_willOverflow : std_logic;
  signal ptrMatch : std_logic;
  signal risingOccupancy : std_logic;
  signal empty : std_logic;
  signal full : std_logic;
  signal pushing : std_logic;
  signal popping : std_logic;
  signal when_Stream_l1011 : std_logic;
  signal when_Stream_l1024 : std_logic;
  signal ptrDif : unsigned(1 downto 0);
begin
  io_push_ready <= io_push_ready_read_buffer;
  io_pop_valid <= io_pop_valid_read_buffer;
  process(pushing)
  begin
    pushPtr_willIncrement <= pkg_toStdLogic(false);
    if pushing = '1' then
      pushPtr_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_flush)
  begin
    pushPtr_willClear <= pkg_toStdLogic(false);
    if io_flush = '1' then
      pushPtr_willClear <= pkg_toStdLogic(true);
    end if;
  end process;

  pushPtr_willOverflowIfInc <= pkg_toStdLogic(pushPtr_value = pkg_unsigned("11"));
  pushPtr_willOverflow <= (pushPtr_willOverflowIfInc and pushPtr_willIncrement);
  process(pushPtr_value,pushPtr_willIncrement,pushPtr_willClear)
  begin
    pushPtr_valueNext <= (pushPtr_value + pkg_resize(unsigned(pkg_toStdLogicVector(pushPtr_willIncrement)),2));
    if pushPtr_willClear = '1' then
      pushPtr_valueNext <= pkg_unsigned("00");
    end if;
  end process;

  process(popping)
  begin
    popPtr_willIncrement <= pkg_toStdLogic(false);
    if popping = '1' then
      popPtr_willIncrement <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_flush)
  begin
    popPtr_willClear <= pkg_toStdLogic(false);
    if io_flush = '1' then
      popPtr_willClear <= pkg_toStdLogic(true);
    end if;
  end process;

  popPtr_willOverflowIfInc <= pkg_toStdLogic(popPtr_value = pkg_unsigned("11"));
  popPtr_willOverflow <= (popPtr_willOverflowIfInc and popPtr_willIncrement);
  process(popPtr_value,popPtr_willIncrement,popPtr_willClear)
  begin
    popPtr_valueNext <= (popPtr_value + pkg_resize(unsigned(pkg_toStdLogicVector(popPtr_willIncrement)),2));
    if popPtr_willClear = '1' then
      popPtr_valueNext <= pkg_unsigned("00");
    end if;
  end process;

  ptrMatch <= pkg_toStdLogic(pushPtr_value = popPtr_value);
  empty <= (ptrMatch and (not risingOccupancy));
  full <= (ptrMatch and risingOccupancy);
  pushing <= (io_push_valid and io_push_ready_read_buffer);
  popping <= (io_pop_valid_read_buffer and io_pop_ready);
  io_push_ready_read_buffer <= (not full);
  when_Stream_l1011 <= (not empty);
  process(when_Stream_l1011,io_push_valid)
  begin
    if when_Stream_l1011 = '1' then
      io_pop_valid_read_buffer <= pkg_toStdLogic(true);
    else
      io_pop_valid_read_buffer <= io_push_valid;
    end if;
  end process;

  when_Stream_l1024 <= pkg_toStdLogic(pushing /= popping);
  ptrDif <= (pushPtr_value - popPtr_value);
  io_occupancy <= unsigned(pkg_cat(pkg_toStdLogicVector((risingOccupancy and ptrMatch)),std_logic_vector(ptrDif)));
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      pushPtr_value <= pkg_unsigned("00");
      popPtr_value <= pkg_unsigned("00");
      risingOccupancy <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      if when_Stream_l1024 = '1' then
        risingOccupancy <= pushing;
      end if;
      if io_flush = '1' then
        risingOccupancy <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamArbiter_1 is
  port(
    io_inputs_0_valid : in std_logic;
    io_inputs_0_ready : out std_logic;
    io_inputs_0_payload_addr : in unsigned(19 downto 0);
    io_inputs_0_payload_id : in unsigned(3 downto 0);
    io_inputs_0_payload_len : in unsigned(7 downto 0);
    io_inputs_0_payload_size : in unsigned(2 downto 0);
    io_inputs_0_payload_burst : in std_logic_vector(1 downto 0);
    io_inputs_0_payload_write : in std_logic;
    io_output_valid : out std_logic;
    io_output_ready : in std_logic;
    io_output_payload_addr : out unsigned(19 downto 0);
    io_output_payload_id : out unsigned(3 downto 0);
    io_output_payload_len : out unsigned(7 downto 0);
    io_output_payload_size : out unsigned(2 downto 0);
    io_output_payload_burst : out std_logic_vector(1 downto 0);
    io_output_payload_write : out std_logic;
    io_chosenOH : out std_logic_vector(0 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamArbiter_1;

architecture arch of StreamArbiter_1 is
  signal io_output_valid_read_buffer : std_logic;

  signal locked : std_logic;
  signal maskProposal_0 : std_logic;
  signal maskLocked_0 : std_logic;
  signal maskRouted_0 : std_logic;
  signal zz_maskProposal_0 : unsigned(0 downto 0);
  signal zz_maskProposal_0_1 : unsigned(1 downto 0);
  signal zz_maskProposal_0_2 : unsigned(1 downto 0);
  signal io_output_fire : std_logic;
begin
  io_output_valid <= io_output_valid_read_buffer;
  maskRouted_0 <= pkg_mux(locked,maskLocked_0,maskProposal_0);
  zz_maskProposal_0 <= unsigned(pkg_toStdLogicVector(io_inputs_0_valid));
  zz_maskProposal_0_1 <= unsigned(pkg_cat(std_logic_vector(zz_maskProposal_0),std_logic_vector(zz_maskProposal_0)));
  zz_maskProposal_0_2 <= (zz_maskProposal_0_1 and pkg_not((zz_maskProposal_0_1 - pkg_resize(unsigned(pkg_toStdLogicVector(maskLocked_0)),2))));
  maskProposal_0 <= pkg_extract(std_logic_vector((pkg_extract(zz_maskProposal_0_2,1,1) or pkg_extract(zz_maskProposal_0_2,0,0))),0);
  io_output_fire <= (io_output_valid_read_buffer and io_output_ready);
  io_output_valid_read_buffer <= (io_inputs_0_valid and maskRouted_0);
  io_output_payload_addr <= io_inputs_0_payload_addr;
  io_output_payload_id <= io_inputs_0_payload_id;
  io_output_payload_len <= io_inputs_0_payload_len;
  io_output_payload_size <= io_inputs_0_payload_size;
  io_output_payload_burst <= io_inputs_0_payload_burst;
  io_output_payload_write <= io_inputs_0_payload_write;
  io_inputs_0_ready <= (maskRouted_0 and io_output_ready);
  io_chosenOH <= pkg_toStdLogicVector(maskRouted_0);
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      locked <= pkg_toStdLogic(false);
      maskLocked_0 <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      if io_output_valid_read_buffer = '1' then
        maskLocked_0 <= maskRouted_0;
      end if;
      if io_output_valid_read_buffer = '1' then
        locked <= pkg_toStdLogic(true);
      end if;
      if io_output_fire = '1' then
        locked <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamFork_1 is
  port(
    io_input_valid : in std_logic;
    io_input_ready : out std_logic;
    io_input_payload_addr : in unsigned(19 downto 0);
    io_input_payload_id : in unsigned(3 downto 0);
    io_input_payload_len : in unsigned(7 downto 0);
    io_input_payload_size : in unsigned(2 downto 0);
    io_input_payload_burst : in std_logic_vector(1 downto 0);
    io_input_payload_write : in std_logic;
    io_outputs_0_valid : out std_logic;
    io_outputs_0_ready : in std_logic;
    io_outputs_0_payload_addr : out unsigned(19 downto 0);
    io_outputs_0_payload_id : out unsigned(3 downto 0);
    io_outputs_0_payload_len : out unsigned(7 downto 0);
    io_outputs_0_payload_size : out unsigned(2 downto 0);
    io_outputs_0_payload_burst : out std_logic_vector(1 downto 0);
    io_outputs_0_payload_write : out std_logic;
    io_outputs_1_valid : out std_logic;
    io_outputs_1_ready : in std_logic;
    io_outputs_1_payload_addr : out unsigned(19 downto 0);
    io_outputs_1_payload_id : out unsigned(3 downto 0);
    io_outputs_1_payload_len : out unsigned(7 downto 0);
    io_outputs_1_payload_size : out unsigned(2 downto 0);
    io_outputs_1_payload_burst : out std_logic_vector(1 downto 0);
    io_outputs_1_payload_write : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamFork_1;

architecture arch of StreamFork_1 is
  signal io_outputs_0_valid_read_buffer : std_logic;
  signal io_outputs_1_valid_read_buffer : std_logic;
  signal io_input_ready_read_buffer : std_logic;

  signal zz_io_outputs_0_valid : std_logic;
  signal zz_io_outputs_1_valid : std_logic;
  signal when_Stream_l817 : std_logic;
  signal when_Stream_l817_1 : std_logic;
  signal io_outputs_0_fire : std_logic;
  signal io_outputs_1_fire : std_logic;
begin
  io_outputs_0_valid <= io_outputs_0_valid_read_buffer;
  io_outputs_1_valid <= io_outputs_1_valid_read_buffer;
  io_input_ready <= io_input_ready_read_buffer;
  process(when_Stream_l817,when_Stream_l817_1)
  begin
    io_input_ready_read_buffer <= pkg_toStdLogic(true);
    if when_Stream_l817 = '1' then
      io_input_ready_read_buffer <= pkg_toStdLogic(false);
    end if;
    if when_Stream_l817_1 = '1' then
      io_input_ready_read_buffer <= pkg_toStdLogic(false);
    end if;
  end process;

  when_Stream_l817 <= ((not io_outputs_0_ready) and zz_io_outputs_0_valid);
  when_Stream_l817_1 <= ((not io_outputs_1_ready) and zz_io_outputs_1_valid);
  io_outputs_0_valid_read_buffer <= (io_input_valid and zz_io_outputs_0_valid);
  io_outputs_0_payload_addr <= io_input_payload_addr;
  io_outputs_0_payload_id <= io_input_payload_id;
  io_outputs_0_payload_len <= io_input_payload_len;
  io_outputs_0_payload_size <= io_input_payload_size;
  io_outputs_0_payload_burst <= io_input_payload_burst;
  io_outputs_0_payload_write <= io_input_payload_write;
  io_outputs_0_fire <= (io_outputs_0_valid_read_buffer and io_outputs_0_ready);
  io_outputs_1_valid_read_buffer <= (io_input_valid and zz_io_outputs_1_valid);
  io_outputs_1_payload_addr <= io_input_payload_addr;
  io_outputs_1_payload_id <= io_input_payload_id;
  io_outputs_1_payload_len <= io_input_payload_len;
  io_outputs_1_payload_size <= io_input_payload_size;
  io_outputs_1_payload_burst <= io_input_payload_burst;
  io_outputs_1_payload_write <= io_input_payload_write;
  io_outputs_1_fire <= (io_outputs_1_valid_read_buffer and io_outputs_1_ready);
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      zz_io_outputs_0_valid <= pkg_toStdLogic(true);
      zz_io_outputs_1_valid <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      if io_outputs_0_fire = '1' then
        zz_io_outputs_0_valid <= pkg_toStdLogic(false);
      end if;
      if io_outputs_1_fire = '1' then
        zz_io_outputs_1_valid <= pkg_toStdLogic(false);
      end if;
      if io_input_ready_read_buffer = '1' then
        zz_io_outputs_0_valid <= pkg_toStdLogic(true);
        zz_io_outputs_1_valid <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

end arch;


--StreamFifoLowLatency_1 replaced by StreamFifoLowLatency

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity BufferCC_3 is
  port(
    io_dataIn : in std_logic;
    io_dataOut : out std_logic;
    io_mainClk : in std_logic
  );
end BufferCC_3;

architecture arch of BufferCC_3 is
  attribute async_reg : string;

  signal buffers_0 : std_logic;
  attribute async_reg of buffers_0 : signal is "true";
  signal buffers_1 : std_logic;
  attribute async_reg of buffers_1 : signal is "true";
begin
  io_dataOut <= buffers_1;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4SharedOnChipRam is
  port(
    io_axi_arw_valid : in std_logic;
    io_axi_arw_ready : out std_logic;
    io_axi_arw_payload_addr : in unsigned(14 downto 0);
    io_axi_arw_payload_id : in unsigned(3 downto 0);
    io_axi_arw_payload_len : in unsigned(7 downto 0);
    io_axi_arw_payload_size : in unsigned(2 downto 0);
    io_axi_arw_payload_burst : in std_logic_vector(1 downto 0);
    io_axi_arw_payload_write : in std_logic;
    io_axi_w_valid : in std_logic;
    io_axi_w_ready : out std_logic;
    io_axi_w_payload_data : in std_logic_vector(31 downto 0);
    io_axi_w_payload_strb : in std_logic_vector(3 downto 0);
    io_axi_w_payload_last : in std_logic;
    io_axi_b_valid : out std_logic;
    io_axi_b_ready : in std_logic;
    io_axi_b_payload_id : out unsigned(3 downto 0);
    io_axi_b_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_valid : out std_logic;
    io_axi_r_ready : in std_logic;
    io_axi_r_payload_data : out std_logic_vector(31 downto 0);
    io_axi_r_payload_id : out unsigned(3 downto 0);
    io_axi_r_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_payload_last : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4SharedOnChipRam;

architecture arch of Axi4SharedOnChipRam is
  signal zz_ram_port0 : std_logic_vector(31 downto 0);
  signal zz_Axi4Incr_result : unsigned(11 downto 0);
  signal zz_Axi4Incr_result_1 : unsigned(10 downto 0);
  signal zz_Axi4Incr_result_2 : unsigned(0 downto 0);
  signal zz_Axi4Incr_result_3 : unsigned(9 downto 0);
  signal zz_Axi4Incr_result_4 : unsigned(1 downto 0);
  signal zz_Axi4Incr_result_5 : unsigned(8 downto 0);
  signal zz_Axi4Incr_result_6 : unsigned(2 downto 0);
  signal zz_Axi4Incr_result_7 : unsigned(7 downto 0);
  signal zz_Axi4Incr_result_8 : unsigned(3 downto 0);
  signal zz_Axi4Incr_result_9 : unsigned(6 downto 0);
  signal zz_Axi4Incr_result_10 : unsigned(4 downto 0);
  signal zz_Axi4Incr_result_11 : unsigned(5 downto 0);
  signal zz_Axi4Incr_result_12 : unsigned(5 downto 0);

  signal unburstify_result_valid : std_logic;
  signal unburstify_result_ready : std_logic;
  signal unburstify_result_payload_last : std_logic;
  signal unburstify_result_payload_fragment_addr : unsigned(14 downto 0);
  signal unburstify_result_payload_fragment_id : unsigned(3 downto 0);
  signal unburstify_result_payload_fragment_size : unsigned(2 downto 0);
  signal unburstify_result_payload_fragment_burst : std_logic_vector(1 downto 0);
  signal unburstify_result_payload_fragment_write : std_logic;
  signal unburstify_doResult : std_logic;
  signal unburstify_buffer_valid : std_logic;
  signal unburstify_buffer_len : unsigned(7 downto 0);
  signal unburstify_buffer_beat : unsigned(7 downto 0);
  signal unburstify_buffer_transaction_addr : unsigned(14 downto 0);
  signal unburstify_buffer_transaction_id : unsigned(3 downto 0);
  signal unburstify_buffer_transaction_size : unsigned(2 downto 0);
  signal unburstify_buffer_transaction_burst : std_logic_vector(1 downto 0);
  signal unburstify_buffer_transaction_write : std_logic;
  signal unburstify_buffer_last : std_logic;
  signal Axi4Incr_validSize : unsigned(1 downto 0);
  signal Axi4Incr_result : unsigned(14 downto 0);
  signal Axi4Incr_highCat : unsigned(2 downto 0);
  signal Axi4Incr_sizeValue : unsigned(2 downto 0);
  signal Axi4Incr_alignMask : unsigned(11 downto 0);
  signal Axi4Incr_base : unsigned(11 downto 0);
  signal Axi4Incr_baseIncr : unsigned(11 downto 0);
  signal zz_Axi4Incr_wrapCase : unsigned(1 downto 0);
  signal Axi4Incr_wrapCase : unsigned(2 downto 0);
  signal when_Axi4Channel_l181 : std_logic;
  signal zz_unburstify_result_ready : std_logic;
  signal stage0_valid : std_logic;
  signal stage0_ready : std_logic;
  signal stage0_payload_last : std_logic;
  signal stage0_payload_fragment_addr : unsigned(14 downto 0);
  signal stage0_payload_fragment_id : unsigned(3 downto 0);
  signal stage0_payload_fragment_size : unsigned(2 downto 0);
  signal stage0_payload_fragment_burst : std_logic_vector(1 downto 0);
  signal stage0_payload_fragment_write : std_logic;
  signal zz_io_axi_r_payload_data : unsigned(12 downto 0);
  signal stage0_fire : std_logic;
  signal zz_io_axi_r_payload_data_1 : std_logic_vector(31 downto 0);
  signal stage1_valid : std_logic;
  signal stage1_ready : std_logic;
  signal stage1_payload_last : std_logic;
  signal stage1_payload_fragment_addr : unsigned(14 downto 0);
  signal stage1_payload_fragment_id : unsigned(3 downto 0);
  signal stage1_payload_fragment_size : unsigned(2 downto 0);
  signal stage1_payload_fragment_burst : std_logic_vector(1 downto 0);
  signal stage1_payload_fragment_write : std_logic;
  signal stage0_rValid : std_logic;
  signal stage0_rData_last : std_logic;
  signal stage0_rData_fragment_addr : unsigned(14 downto 0);
  signal stage0_rData_fragment_id : unsigned(3 downto 0);
  signal stage0_rData_fragment_size : unsigned(2 downto 0);
  signal stage0_rData_fragment_burst : std_logic_vector(1 downto 0);
  signal stage0_rData_fragment_write : std_logic;
  signal when_Stream_l342 : std_logic;
  type ram_type is array (0 to 8191) of std_logic_vector(7 downto 0);
  signal ram_symbol0 : ram_type := (
     "00110111","00010011","11100111","00010011","00000000","00000000","00000000","00000000","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00010011","11101111","10000011","10000011","00000011","10000011","00000011","10000011",
     "00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00010011","01110011","10010111","10010011","00010111","00010011",
     "00010111","00010011","10010011","01100011","00100011","00010011","01101111","00010111","00010011","00010011","10010111","10010011","01100011","10000011","00010011","00100011",
     "11100111","00000011","01101111","00010011","00110111","00010011","01110011","00110111","00010011","01110011","11101111","01101111","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00011000","11110100","11111100","00000100","00010000","11101000","10101100","00110100","00110100","10100000","00110100","00110100","00110100","00110100","00110100","00110100",
     "00110100","10010100","00110100","10001000","00110100","00110100","00011000","11010100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100",
     "00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","00101100","01101000","00101100",
     "00101100","00101100","00101100","00101100","00101100","00101100","00101100","01011100","00101100","11100100","10111000","00101100","00101100","00101100","00101100","10111000",
     "00101100","00101100","00101100","00101100","00101100","11011000","10111100","00101100","00101100","10101000","00101100","10011100","00101100","00101100","01010000","11010100",
     "00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100",
     "00110100","00110100","00110100","00110100","00110100","00110100","01101100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00110100","00111000",
     "00110100","11101000","10111100","00110100","00110100","00110100","00110100","10111100","00110100","00110100","00110100","00110100","00110100","11011100","11000000","00110100",
     "00110100","10101100","00110100","10100000","00110100","00110100","01110000","00110000","00110100","00111000","01100011","01100111","01101011","01101111","01110011","01110111",
     "00000000","00110000","00110100","00111000","01000011","01000111","01001011","01001111","01010011","01010111","00000000","00111100","01001100","01110110","01101001","00111010",
     "01101111","01110011","01110010","01101001","01100001","01110101","00001010","01110110","01101001","00111010","01100101","01101001","01100011","01101101","00100000","00100000",
     "01110010","01101111","00101110","01101001","01100001","01100001","01110011","00100000","01100101","00001010","00001010","01010010","00111010","01101100","01110000","01100101",
     "01110101","01110010","01101110","01110011","00100000","00100000","01100101","00100000","01110100","00000000","01010011","01110100","01101101","00000000","00110110","01100101",
     "01110010","01100011","01110101","01100001","01100101","01110011","01110010","01110010","01110010","00000000","00110110","01100001","01100001","01101110","01101110","01110010",
     "01110100","00100000","00100000","01100101","01101011","01010000","01101001","01100111","01110010","01101111","01110101","01100001","01100101","01110011","01110010","01110010",
     "01110010","00000000","00110010","01100101","01110010","01100011","01110101","01100001","01100101","01110011","01110010","01110010","01110010","00000000","00110010","01100001",
     "01100001","01101110","01101110","01110010","01110100","00100000","00100000","01100101","01101011","01011011","01000101","01010010","01101001","01100011","00110000","00110100",
     "00100000","01110101","01100010","01111000","01111000","01011011","01000101","01010010","01100001","01111000","01100011","00100101","00100000","01101000","01100100","00100000",
     "00110000","00000000","01011011","01000101","01010010","01110100","00100000","00100000","00110000","00101101","01101111","00100000","00110000","00110100","01000011","01001101",
     "00100000","01100101","00100000","01101100","01010100","01101100","01100011","00100000","00100000","01101100","01010100","01101100","01101101","01110011","00101001","01100100",
     "01001001","01100001","01101110","01100101","00100000","01100100","01000101","01010010","01110101","01100101","01110101","01100110","01100001","01100101","00100000","01110011",
     "00100000","00100000","01100001","00100000","01110101","00001010","01001001","01100001","01101110","00100000","00100000","01101100","01000111","00101110","00000000","01000011",
     "01101001","00100000","01110011","00100000","01110011","00101101","01100101","01101100","01110011","01101101","01100110","00000000","01000011","01101001","00100000","01100111",
     "00100000","01110011","01010011","01001011","01001101","01110010","01101111","01101001","00100000","01110011","01110011","01100011","00100000","00100000","00100000","01111000",
     "01111000","01011011","01100011","01101001","00100000","00100000","00110000","00110100","01011011","01100011","01100001","01111000","00100000","00110000","00110100","01011011",
     "01100011","01110100","00100000","00100000","00110000","00110100","01011011","01100011","01101001","00100000","00100000","00110000","00110100","01000011","01100101","01101111",
     "01100001","01101110","01101100","01110100","00100000","00100000","01000100","01101101","01101111","01110101","01101110","01100101","01110100","00100000","01100101","00000000",
     "01000101","01110010","01100101","01110100","00000000","01000011","01101111","01100001","01100001","01101111","01100001","01101110","01110010","01100101","01110011","00100000",
     "01110101","00100000","01100001","01100011","01100001","01110111","00100000","01110101","00100000","01100001","01101111","01110000","01100110","00101110","01010011","01101001",
     "01001000","00000000","01010011","01101011","01001000","01001000","11111000","11111000","00011100","01110100","01111100","10000100","10001100","01000100","01010000","01011100",
     "01101000","00010100","00100000","00101100","00111000","11100100","11110000","11111100","00001000","01010100","01100101","00000000","00101101","00101011","00000000","00110001",
     "00110100","00000000","00110011","01100101","00000000","00110101","00110000","00000000","00101101","00110011","00000000","00101101","00101011","00000000","00101011","01100101",
     "00000000","00110011","00110100","00000000","00101110","00110100","00000000","00101101","00101110","00000000","00101011","00110100","00000000","00110101","00000000","00110001",
     "00000000","00101101","00000000","00101011","00000000","00000000","00000011","00000100","00000100","00000101","00000101","00000101","00000101","00000110","00000110","00000110",
     "00000110","00000110","00000110","00000110","00000110","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",
     "00000111","00000111","00000111","00000111","00000111","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00000000","00000001","01100110","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","10010011","01100011","10110111","10010011","00010011","00110011","10000011","01100111","10110111","00000011","01100111","00000011","01100111","00000011",
     "01100111","10110111","00000011","01100111","00000011","01100111","00010011","01100111","10110011","10010011","00010011","10010011","01100011","10110111","10010011","10110011",
     "10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","10110011","10010011","00010011","10010011",
     "01100011","10110111","10010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011",
     "10110011","10010011","00010011","10010011","01100011","10110111","10010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111",
     "00010011","10110011","10010011","10010011","10110011","10010011","00010011","10010011","01100011","10110111","10010011","10110011","10010011","10010011","10010011","00010011",
     "01100011","10110111","10010011","10110011","00010011","00010011","01100111","00110011","10010011","00010011","00010011","10010011","01100011","00110111","00010011","10110011",
     "10010011","10010011","00110011","00010011","10010011","00010011","01100011","00110111","00010011","10110011","10010011","10010011","00110011","00010011","00010011","10010011",
     "01100011","00110111","00010011","10110011","10010011","10010011","00110011","00010011","00010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011",
     "00110011","00010011","00010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","00110011","00010011","00010011","10010011","01100011","00110111",
     "00010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","00010011","10010011",
     "01100011","00110111","00010011","10110011","10010011","10010011","00010011","00110011","00010011","00010011","10010011","00010011","01100011","10110111","10010011","00110011",
     "00010011","00010011","10110011","10010011","10010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","10110011","10010011","10010011","00010011",
     "01100011","10110111","10010011","00110011","00010011","00010011","10110011","10010011","10010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011",
     "10110011","10010011","10010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","10110011","10010011","10010011","00010011","01100011","10110111",
     "10010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","10010011","00010011",
     "01100011","10110111","10010011","00110011","00010011","00010011","01100111","00110011","10010011","00010011","00010011","00010011","00010011","10010011","01100011","10110111",
     "10010011","10110011","10010011","10010011","00110011","10010011","10010011","00010011","01100011","10110111","10010011","10110011","10010011","10010011","00110011","00010011",
     "10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","10110011","10010011","00010011","10010011","01100011","10110111","10010011","10110011",
     "10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","10110011","10010011","00010011","10010011",
     "01100011","10110111","10010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011",
     "00010011","10010011","01100011","10110111","10010011","10110011","10010011","10010011","00010011","10110011","10010011","00010011","00010011","10010011","01100011","10110111",
     "10010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","10110011","10010011",
     "00010011","10010011","01100011","10110111","10010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011","01100011","00110111","00010011","10110011",
     "10010011","10010011","10110011","10010011","00010011","10010011","01100011","10110111","10010011","10110011","10010011","10010011","00110011","00010011","10010011","10010011",
     "01100011","00110111","00010011","10110011","10010011","10010011","10110011","10010011","00010011","10010011","01100011","10110111","10010011","10110011","10010011","10010011",
     "10010011","10010011","01100011","00110111","00010011","10110011","10010011","10010011","00010011","10110011","00010011","10010011","10010011","10010011","00010011","00010011",
     "01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011",
     "10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111",
     "00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011",
     "10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011",
     "00010011","00010011","10010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","10010011","00110011","00010011","10010011","10010011","00010011",
     "01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011",
     "00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111",
     "10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011",
     "00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011",
     "00010011","00010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","01100111","00110011","00010011","10010011","00010011","10010011",
     "10010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","10110011","00010011","00010011","10010011","01100011","10110111","10010011","00110011",
     "00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011",
     "01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011",
     "00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111",
     "10010011","00110011","00010011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10010011","00110011","00010011","10010011",
     "10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011",
     "00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011","10110011","10010011","00010011","00010011",
     "01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111","00010011","00110011","00010011","00010011",
     "10110011","10010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","00110011","00010011","10010011","00010011","01100011","00110111",
     "00010011","00110011","00010011","00010011","00010011","00010011","01100011","10110111","10010011","00110011","00010011","00010011","01100111","00010011","01100111","00010011",
     "00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00010011","10010011","00010011",
     "01100011","10110111","10010011","00010011","01100011","00010011","00010011","00010011","01100011","00010011","10010011","01100011","01100011","00010011","01100011","10010011",
     "00010011","01100011","10010011","00010011","01100011","10010011","01100011","10010011","10010011","10110011","01100011","10010011","00100011","00010011","10010011","10010011",
     "00010011","10010011","01100011","10010011","00110011","10010011","01100011","01100011","00010011","00010011","10010011","00100011","11101111","00000011","10110011","10010011",
     "00010011","01100011","00100011","10010011","01100011","10010011","01100011","10010011","01100011","01100011","01100011","00010011","00010011","00110011","00010011","00010011",
     "00010011","00010011","10010011","00110011","11101111","10110011","10010011","01100011","10110011","00010011","00010011","10010011","11101111","10110011","00110011","00010011",
     "00010011","00010011","10000011","10110011","10110011","10100011","10110011","00010011","11100011","10110011","01100011","10010011","10010011","00110011","00010011","00010011",
     "00010011","10010011","11101111","10110011","10000011","00000011","00010011","00000011","10000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011",
     "00000011","10000011","00010011","01100111","10010011","00010011","00010011","00010011","10010011","01100011","01101111","10110111","10010011","01101111","00010011","01101111",
     "10110011","10010011","00010011","11100011","00010011","00010011","01101111","00010011","10110011","10010011","00110011","00010011","10010011","10110011","10000011","10110011",
     "10100011","11100011","01101111","10010011","00010011","01101111","10010011","00100011","10010011","10100011","10010011","01101111","10010011","01101111","10010011","00100011",
     "10010011","01101111","00010011","10010011","01101111","10010011","00010011","10010011","01101111","10010011","01100011","00110111","10000011","10010011","10010011","11100011",
     "00100011","01100111","00110111","10000011","10010011","10010011","11100011","10010011","00100011","01101111","00010011","00100011","00100011","00100011","00100011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","10000011",
     "00010011","00100011","11100011","00010011","10110111","00110111","10110111","00010011","00010011","10010011","00010011","10010011","10110111","00010011","01100011","00100011",
     "10000011","00010011","00010011","11100011","00100011","10000011","01100011","00010011","10010011","00110111","00010011","00110011","01100011","10000011","10010011","10010011",
     "11100011","00110011","00100011","00010011","10000011","11100011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011",
     "10000011","00000011","10000011","00010011","01100111","10000011","10010011","10010011","11100011","00100011","01101111","10000011","10010011","10010011","00010011","00010011",
     "10010011","01100011","00010011","00110011","00000011","01100111","10010011","00010011","10000011","10010011","00010011","00010011","11100011","00010011","00010011","10010011",
     "01100011","00010011","10010011","01100011","00010011","00010011","01100011","00010011","00010011","01100011","00010011","00010011","00010011","01100011","00010011","00110011",
     "00000011","01100111","10010011","00010011","01101111","10010011","00010011","01101111","10010011","00010011","01101111","10010011","00010011","01101111","00000011","00010011",
     "10010011","00010011","00010011","01100011","00110111","00010011","00010011","00110011","00000011","01100111","10000011","00010011","00010011","00010011","00010011","01100011",
     "00010011","01100011","10010011","00010011","01101111","10010011","00010011","00010011","10110011","10010011","10010011","10110011","10000011","10010011","00010011","00010011",
     "11100011","01101111","10000011","10010011","10000011","00010011","11100011","10110011","10010011","01101111","10010011","10010011","00010011","00010011","10000011","00010011",
     "00010011","11101111","10000011","00010011","00010011","11100011","01101111","10010011","00010011","01101111","10010011","00000011","00010011","01100011","00000011","11100011",
     "11100011","00010011","01101111","10110011","01100011","00010011","10000011","11100011","10010011","10110011","01100011","01100011","00010011","00010011","00110011","00110011",
     "10010011","00010011","00010011","10010011","00110011","10010011","10110011","11100011","10110011","10010011","11100011","10010011","10010011","00010011","10110011","00000011",
     "00010011","10010011","00100011","11100011","10010011","00110011","00110011","00110011","01100011","00000011","10010011","00100011","01100011","10000011","10010011","10100011",
     "01100011","10000011","00100011","00010011","00010011","01100011","10110011","00010011","00010011","10010011","11101111","00110011","10000011","11100011","01101111","10010011",
     "00010011","01100011","10000011","00010011","00010011","01101111","10010011","00010011","01101111","10010011","10010011","10010011","01100011","10000011","00010011","00010011",
     "00100011","00010011","01100011","00010011","10010011","00010011","11101111","10000011","00110011","11100011","01101111","00010011","10010011","10010011","00010011","01100011",
     "00100011","00000011","01100011","00010011","00100011","10000011","11100011","00010011","01101111","00010011","00010011","00010011","00110011","00010011","00010011","00110011",
     "10000011","00010011","00010011","00010011","11100011","10010011","01101111","00000011","10000011","00010011","00010011","00010011","00110011","10010011","01101111","00010011",
     "10010011","00010011","00010011","11100011","01101111","00010011","00000011","10010011","00010011","01100011","00110111","00010011","00000011","00000011","00000011","00000011",
     "10000011","10000011","10010011","10010011","10010011","00010011","10010011","00010011","00010011","00010011","00010011","10010011","00010011","00110011","00110011","10110011",
     "10110011","10110011","00110011","00110011","00110011","10110011","10110011","00000011","10000011","10000011","10000011","10000011","00000011","00000011","00000011","10000011",
     "00000011","00110011","00000011","00010011","10010011","10100011","00100011","10100011","00100011","10100011","00100011","00100011","10100011","00100011","00100011","10100011",
     "10100011","00100011","00100011","10100011","00110011","10100011","00000011","10010011","00010011","00100011","01100011","10010011","01100011","00010011","00010011","10010011",
     "00010011","00100011","11101111","00010011","10010011","00110011","11101111","10000011","00110011","10000011","00010011","00010011","11100011","01101111","00010011","00000011",
     "00010011","01100011","00010011","01101111","10010011","00010011","01101111","00000011","00010011","00000011","01100011","10010011","01100011","00010011","10110011","00010011",
     "10010011","00010011","00010011","00110011","00110011","00110011","00000011","00100011","00110011","00000011","00110011","10100011","00110011","00000011","00010011","00110011",
     "00100011","00010011","00000011","00110011","00010011","00100011","01100011","00010011","01100011","00010011","10010011","00010011","00110011","10010011","00110011","00110011",
     "00110011","00110011","00000011","00100011","00110011","00000011","00110011","00100011","00110011","00000011","00010011","00110011","00010011","00100011","10010011","00000011",
     "00110011","10010011","00100011","10010011","01100011","00010011","01100011","00010011","10010011","00010011","00110011","10010011","00110011","00110011","00110011","00110011",
     "00000011","00100011","00110011","00000011","00110011","00100011","00110011","00000011","00010011","00110011","00010011","00100011","00000011","00010011","10110011","00010011",
     "00100011","00010011","01100011","00010011","01100011","00010011","00010011","00010011","00110011","00010011","10110011","00110011","00110011","00110011","00000011","00100011",
     "00110011","00000011","00110011","00100011","00110011","10000011","00010011","00110011","00010011","00100011","10010011","10010011","01100011","01100011","00110011","00010011",
     "00010011","10010011","00100011","11101111","10000011","00110011","10110011","10110011","10010011","00010011","00010011","10010011","00100011","11101111","10000011","00110011",
     "00010011","01100011","00010011","10010011","00010011","10110011","10110011","10100011","10110011","11100011","10000011","00010011","01100011","01101111","10010011","00010011",
     "10010011","10000011","00010011","00010011","01101111","00000011","10010011","00010011","01101111","10010011","00010011","00010011","00100011","10000011","00010011","00010011",
     "01100011","01101111","10010011","10010011","01101111","01100011","00010011","00010011","10010011","00110011","11101111","10010011","01101111","00010011","01101111","00010011",
     "01100011","10110011","00010011","00010011","10010011","00100011","11101111","10000011","00110011","10110011","10110011","01101111","00010011","00100011","00010011","00010011",
     "00000011","00110011","00010011","00100011","10010011","11100011","00010011","00110011","10010011","00100011","00010011","10010011","00000011","00110011","10010011","00100011",
     "10010011","11100011","00010011","00110011","10010011","00100011","00010011","00010011","00000011","10110011","00010011","00100011","00010011","11100011","00010011","00110011",
     "00010011","00010011","00100011","01101111","10010011","10010011","00010011","00010011","10010011","00010011","00100011","11101111","10000011","10010011","00010011","11100011",
     "10010011","00010011","10010011","00010011","10110011","10110011","10100011","10110011","11100011","01101111","00010011","00010011","01101111","10010011","01101111","00010011",
     "11100011","00010011","00110011","10010011","10110011","10010011","00110011","00000011","00110011","00100011","01101111","00010011","11100011","00010011","00110011","10010011",
     "10110011","10010011","00110011","00000011","00110011","00100011","01101111","10010011","11100011","00010011","10110011","00010011","00110011","00010011","10110011","10000011",
     "00110011","00100011","01101111","10010011","01100011","00010011","00110011","10010011","00010011","00010011","00110011","00000011","00110011","00100011","01101111","10010011",
     "00010011","00010011","01101111","10010011","11100011","10010011","01101111","10000011","00010011","00010011","00100011","00010011","10000011","00010011","01100011","01101111",
     "10010011","01101111","00110011","00010011","10000011","00010011","10100011","11100011","01101111","10010011","10010011","10010011","01101111","00010011","00100011","00100011",
     "00100011","00100011","00100011","00000011","10010011","10010011","00010011","01100011","10010011","10010011","10010011","10010011","00010011","10110011","10010011","10000011",
     "01100011","10010011","01100011","00010011","00010011","00010011","10010011","00010011","00010011","11101111","00110011","00100011","00010011","00100011","10000011","00000011",
     "00010011","10000011","00000011","10000011","00010011","01100111","10010011","00010011","01100011","00010011","10000011","00000011","10000011","00000011","00010011","11101111",
     "10000011","00010011","00010011","01100011","00100011","10000011","01101111","00010011","00010011","11101111","10000011","00010011","00010011","11100011","10000011","00100011",
     "01101111","00010011","00100011","00100011","00100011","00100011","00100011","00100011","00000011","00010011","10010011","10010011","10010011","00010011","01100011","10010011",
     "10010011","10010011","00010011","10110011","10010011","10000011","01100011","10010011","01100011","00010011","00010011","00010011","10010011","00010011","00010011","11101111",
     "00110011","00100011","00010011","00100011","00000011","10010011","10010011","10010011","01100011","10010011","10010011","10010011","00010011","10110011","10000011","01100011",
     "10010011","01100011","00010011","00010011","10010011","10010011","10010011","00010011","11101111","00110011","00100011","00010011","00100011","10000011","00000011","00110011",
     "10000011","00000011","10000011","00000011","00010011","01100111","10010011","00010011","01100011","00010011","10000011","00000011","10000011","00000011","00010011","11101111",
     "10000011","00010011","00010011","01100011","00100011","10000011","01101111","10010011","00010011","01100011","00010011","10000011","00000011","10000011","00000011","00010011",
     "11101111","10000011","10010011","10010011","01100011","00100011","10000011","01101111","00010011","00010011","11101111","10000011","00010011","00010011","11100011","10000011",
     "00100011","01101111","00010011","00010011","11101111","10000011","10010011","10010011","11100011","10000011","00100011","01101111","01100011","00000011","10000011","00110011",
     "01100111","10000011","00010011","00010011","00010011","10010011","10110011","00100011","10000011","00010011","00010011","00010011","10010011","10110011","00100011","00000011",
     "10000011","00110011","01100111","10000011","00100011","10000011","00100011","01100111","00010011","00100011","00100011","00100011","00100011","00100011","00100011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00100011","10000011","00100011","00010011","00000011","01100011","00100011","00010011","00010011","00010011","00010011",
     "10000011","10010011","00100011","01100011","01100011","00000011","10010011","10010011","00000011","01100011","01101111","00000011","10000011","00000011","01100011","10000011",
     "11100011","10010011","01101111","10010011","00010011","00000011","00100011","11100011","01100011","00000011","00010011","00010011","00000011","00010011","10010011","01100011",
     "00010011","00010011","00110011","00010011","00010011","10000011","01100011","00000011","00100011","10000011","00100011","00100011","10000011","01100011","00010011","10010011",
     "10010011","00100011","00010011","00010011","00010011","11100011","10010011","10110011","10110011","10010011","10010011","00100011","01100011","10000011","10010011","00000011",
     "00000011","10000011","00100011","00100011","00000011","00000011","00100011","10000011","00100011","01100011","10000011","00000011","10000011","01100011","10000011","11100011",
     "10000011","01100011","10000011","10000011","00000011","11101111","10000011","00100011","11100011","10000011","10000011","00000011","00010011","00100011","10000011","00100011",
     "10010011","00100011","00100011","00010011","10010011","00010011","00010011","10010011","10010011","10000011","10010011","01100011","11100011","10010011","00010011","00010011",
     "00010011","01100011","01100011","01100011","10000011","00000011","10000011","00010011","00010011","00010011","10010011","10110011","00100011","10000011","10000011","00010011",
     "00010011","10010011","00010011","10110011","00100011","10000011","10110011","01100011","10010011","00000011","00010011","01100011","00100011","10010011","11100011","01100011",
     "01100011","10010011","00010011","00000011","11100011","10010011","10010011","01101111","10000011","00000011","10000011","11100011","10000011","11100011","10000011","11100011",
     "01101111","10010011","10010011","00000011","01101111","11100011","00100011","01100011","00010011","01100011","00010011","00010011","10010011","10010011","01101111","01100011",
     "00000011","10010011","00000011","01100011","01101111","00000011","10000011","00000011","11100011","10000011","11100011","01101111","00000011","10010011","00010011","00000011",
     "00010011","00010011","00110011","00010011","00010011","01101111","00000011","01100011","10000011","10000011","00000011","11101111","00000011","00100011","11100011","10000011",
     "00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00010011","01100111","00100011","00100011",
     "11100011","01100011","10010011","00100011","10010011","00100011","00010011","00010011","00010011","00100011","00010011","10000011","10010011","10010011","10010011","00100011",
     "10000011","10010011","01100011","10000011","11100011","10000011","01100011","01100011","01100011","10000011","10000011","10000011","10010011","00010011","01100011","10010011",
     "10010011","10010011","00010011","10110011","10000011","01100011","01100011","00010011","00010011","00010011","10010011","11101111","00010011","10010011","10110011","00100011",
     "10010011","00100011","10000011","10010011","10010011","01100011","10010011","10010011","10010011","00010011","10110011","10000011","01100011","01100011","00010011","00010011",
     "10010011","10010011","11101111","10010011","10010011","10110011","00100011","10010011","00100011","10110011","01100011","10010011","10000011","10010011","01100011","00100011",
     "00010011","11100011","01100011","01100011","10010011","10010011","10000011","11100011","00010011","00010011","01101111","10010011","10010011","00000011","01101111","00010011",
     "11100011","00000011","00100011","10010011","11100011","10000011","10010011","00100011","11100011","00100011","01110011","00000011","00010011","11101111","10000011","10010011",
     "10010011","01100011","10000011","00100011","01101111","10010011","00010011","01100011","00010011","10000011","00000011","10000011","00000011","00010011","11101111","10000011",
     "10010011","10010011","01100011","00100011","10000011","01101111","00000011","00010011","11101111","10000011","00010011","00010011","01100011","10000011","00100011","01101111",
     "10010011","00010011","01100011","00010011","10000011","00000011","10000011","00000011","00010011","11101111","10000011","00010011","00010011","01100011","00100011","10000011",
     "01101111","00000011","01101111","10000011","01110011","10010011","00110011","00100011","10110111","00010011","10010011","10010011","00010011","00010011","00110011","00100011",
     "00100011","00000011","10010011","10110011","00100011","00010011","01100011","00010011","00000011","01100011","00100011","00100011","00100011","00010011","10010011","00100011",
     "00100011","00000011","01100011","10010011","10110111","10010011","10010011","10010011","00010011","01100011","10010011","01100011","00010011","00010011","10110011","10010011",
     "10010011","00010011","00100011","10110011","00100011","00010011","00100011","10110011","00100011","00100011","00000011","00010011","10010011","10010011","11100011","10000011",
     "01100011","10010011","00110011","00110111","10010011","00010011","10000011","01100011","00100011","00000011","10010011","10000011","11100011","10010011","10010011","10010011",
     "10010011","10010011","00010011","00010011","00010011","00010011","00000011","00010011","01100011","11100011","10010011","00010011","10010011","01100011","01100011","01100011",
     "00000011","00000011","00000011","00010011","00010011","00010011","00010011","00110011","00100011","00000011","10000011","10010011","10010011","00010011","10010011","00110011",
     "00100011","00000011","00110011","01100011","00010011","10000011","00010011","01100011","00100011","10010011","11100011","01100011","01100011","00010011","00010011","10000011",
     "11100011","10010011","10010011","01101111","00010011","00010011","10000011","01101111","11100011","00100011","01100011","10010011","11100011","00100011","01110011","00010011",
     "00010011","10010011","10010011","10010011","00110011","10110011","10110011","00100011","00000011","10010011","10000011","11100011","01101111","00010011","01100111","00000011",
     "00010011","10010011","01101111","00010011","10010011","01101111","00000011","10010011","01100011","00000011","00010011","01100011","00100011","10000011","00100011","00100011",
     "10000011","00010011","00100011","10010011","00100011","00000011","10000011","00100011","00000011","00100011","01100111","00010011","00010011","01100111","00000011","10000011",
     "10010011","00000011","00010011","00100011","00100011","10000011","10000011","00100011","00100011","01100111","00000011","10000011","00100011","00000011","00100011","00100011",
     "00100011","01100111","00000011","01100011","01100011","10000011","10000011","01100011","01101111","10000011","10000011","01100011","00000011","11100011","01100111","11100011",
     "10000011","00000011","10000011","01100011","01101111","10000011","10000011","01100011","00000011","11100011","01101111","01100111","01100111","01100111","01100011","00010011",
     "01101111","00010011","10000011","00100011","00010011","11100011","01100111","01100011","00010011","00100011","00100011","00100011","00100011","00100011","00100011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00010011","10010011","00010011","10010011","00010011","00010011","10010011","00010011","00010011","10010011","00010011",
     "10010011","00000011","10010011","01100011","11100011","10010011","01100011","01100011","01100011","10000011","00000011","00010011","11100111","01100011","10010011","00000011",
     "10010011","01100011","00100011","00010011","11100011","01100011","01100011","10010011","10010011","00000011","11100011","00010011","00010011","01101111","10010011","10010011",
     "00000011","01101111","00010011","11100011","00100011","01100011","10010011","11100011","00100011","01110011","10000011","00000011","00010011","10000011","00000011","10000011",
     "00000011","10000011","00000011","10000011","00000011","10000011","00000011","00010011","01100111","00100011","01110011","00010011","10010011","01100111","00110111","10010011",
     "00010011","00100011","00100011","10110111","00100011","10110111","00100011","00110111","10010011","00100011","10010011","00100011","00010011","00100011","01100111","10110111",
     "00000011","10110111","00100011","00100011","01100111","10110111","00110111","10000011","00000011","10000011","00000011","00110011","10110011","10110011","10110011","01100111",
     "00010011","00010011","10010011","00100011","11101111","10000011","00010011","01100111","00010011","00100011","00010011","00110111","10010011","00010011","00100011","11101111",
     "00110111","10010011","00010011","11101111","10010011","00100011","10000011","00000011","00010011","01100111","00100011","00110111","00010011","01101111","01100111","00010011",
     "00100011","00100011","00100011","00100011","00000011","00100011","00100011","00010011","10010011","01100011","10010011","00010011","11101111","10000011","11101111","00100011",
     "10010011","00010011","11101111","10000011","11101111","00100011","01100011","10010011","11100011","10000011","00000011","10000011","00000011","00010011","00010011","01100111",
     "00100011","10010011","11100011","10010011","01101111","10000011","01100011","00110111","10000011","10010011","10010011","11100011","00100011","00010011","10000011","11100011",
     "01100111","10000011","01100011","00110111","10000011","10010011","10010011","11100011","00100011","00010011","10000011","11100011","00110111","10000011","10010011","10010011",
     "11100011","10010011","00100011","01100111","00010011","10010011","00010011","01100011","10010011","10010011","10010011","10010011","10010011","10010011","10110111","10110111",
     "00010011","00010011","10010011","00010011","10010011","10010011","00010011","10010011","00010011","01100011","10010011","10110011","10000011","00010011","00110011","10010011",
     "10010011","01100111","10010011","00000011","10010011","01100011","10010011","10000011","10110011","00100011","00000011","10100011","00000011","00100011","00000011","10100011",
     "01100011","00000011","00100011","00000011","10100011","00000011","00100011","01100011","00000011","10100011","10110011","00100011","10010011","10010011","10010011","00010011",
     "10010011","00010011","00010011","11100011","00010011","10010011","00110011","10010011","10010011","00000011","10010011","01100011","10010011","01101111","10010011","00000011",
     "10010011","11100011","01100011","00110011","10010011","00110011","01101111","10010011","00000011","10010011","11100011","11100011","01100111","00010011","00110011","10010011",
     "00110011","01101111","10000011","10000011","01100011","00010011","00010011","01100011","10000011","00010011","00010011","00010011","10010011","01100011","00100011","10000011",
     "01100011","10010011","01100011","00010011","00010011","10010011","00010011","00010011","01100011","01100011","10000011","00010011","00010011","01100011","01100011","10010011",
     "00010011","00010011","11100011","10000011","10010011","00100011","10000011","01100011","00010011","00010011","01100011","00010011","10010011","00010011","00010011","10010011",
     "00010011","01100011","01100011","10000011","00010011","10010011","10010011","00100011","00100011","00010011","01100111","00010011","01100011","00010011","01100011","00010011",
     "01100011","10000011","00100011","10010011","10010011","00100011","00100011","00010011","01100111","10000011","00010011","10010011","10010011","00100011","00100011","00010011",
     "01100111","00100011","10000011","01100011","00010011","01100011","00000011","10010011","10010011","00010011","00010011","01100011","10010011","01100011","00100011","10010011",
     "00100011","00010011","01100111","00100011","10000011","01100011","00010011","10010011","11100011","00010011","10010011","01101111","00000011","00010011","00100011","10000011",
     "01100011","00010011","00010011","01100011","10000011","10010011","10010011","10010011","00100011","01100011","10010011","00100011","00010011","01100111","10000011","01100011",
     "00010011","01100011","10000011","10010011","10010011","10010011","10010011","00100011","11100011","10000011","01100011","10010011","01100011","00010011","10010011","10010011",
     "10010011","01100011","10000011","00010011","10010011","10010011","00100011","01101111","10000011","00010011","00010011","01100011","01100011","10010011","01101111","10000011",
     "00010011","10010011","01100011","01100011","00010011","01101111","00100011","10000011","01100011","00010011","01100011","10010011","01101111","00100011","10000011","01100011",
     "10010011","00010011","11100011","00010011","10010011","01101111","10010011","01101111","00010011","10010011","01101111","10010011","01101111","00010011","10010011","01101111",
     "00010011","10010011","01101111","10010011","01101111","00010011","10010011","01101111","00010011","10010011","01101111","00010011","10010011","01101111","00010011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00010011","10000011","10010011","00100011","00100011","00100011","00100011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","10010011","00010011","00010011","00010011",
     "10010011","01100011","10010011","10010011","00010011","11101111","10010011","00010011","00110011","00000011","10000011","00000011","10010011","00100011","11100011","00100011",
     "10110011","10000011","01100011","10010011","10010011","00110011","01100011","00100011","10000011","10110011","00100011","01100011","10000011","00110011","11100011","10110011",
     "00100011","11100011","10000011","00100011","10010011","01100011","10010011","00010011","11101111","10010011","00010011","00110011","00000011","10000011","00000011","10010011",
     "00100011","11100011","00100011","01100011","10010011","10000011","00110011","01100011","00100011","00000011","00110011","00100011","11100011","00010011","00010011","00000011",
     "10010011","00010011","11101111","10010011","00000011","00010011","11101111","10010011","11100011","10000011","00000011","10000011","00000011","10000011","00000011","10000011",
     "00000011","10000011","00010011","01100111","00110011","00100011","11100011","01101111","10110011","11100011","01101111","11100011","01101111","00010011","00100011","00100011",
     "10110111","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","10110011","01100011","00010011","10110011","00010011",
     "10010011","10110011","10010011","00010011","10010011","00010011","10010011","10010011","00010011","00010011","10010011","00110011","10010011","10000011","10010011","10110011",
     "00100011","11100011","00010011","00110011","01100011","00010011","01101111","00110011","00010011","10010011","00010011","00010011","00010011","10110011","00010011","10010011",
     "10000011","00010011","10010011","10110011","00100011","11100011","10010011","00110011","10110011","01100011","00010011","01101111","00110011","10010011","00010011","10010011",
     "00010011","10010011","00010011","00110011","10010011","01101111","00010011","10010011","00010011","10010011","01100011","00000011","00010011","00010011","10110011","00110011",
     "10010011","00110011","11100011","00010011","10010011","00010011","00010011","10010011","11100011","10010011","10110011","01100011","10010011","01101111","10010011","11101111",
     "10010011","00010011","00110011","10010011","00100011","10010011","00010011","10010011","00000011","00000011","10010011","00010011","00110011","10110011","00100011","11100011",
     "10010011","00110011","11100011","00010011","00010011","10010011","10010011","00010011","00010011","00010011","01101111","00010011","00010011","00010011","00010011","10010011",
     "01100011","00000011","00010011","00010011","10110011","10110011","10010011","00110011","11100011","00010011","00010011","00010011","10010011","00010011","10010011","11100011",
     "00010011","00110011","11100011","11101111","10010011","10010011","10010011","00010011","00010011","10010011","00010011","00100011","00010011","00010011","10010011","00010011",
     "10000011","00000011","00010011","00010011","10110011","00110011","10110011","00100011","11100011","00010011","10010011","00010011","11100011","00010011","10110011","10110011",
     "11100011","00010011","00010011","10010011","10010011","00010011","00010011","00010011","01101111","00010011","00010011","00010011","00010011","10010011","01100011","00000011",
     "00010011","00010011","10110011","10110011","10010011","00110011","11100011","00010011","00010011","00010011","10010011","00010011","10010011","11100011","00010011","00110011",
     "11100011","11101111","10010011","00010011","10010011","00010011","00010011","00100011","00010011","10010011","00010011","10010011","00000011","10000011","10010011","10010011",
     "10110011","00110011","00010011","10010011","00010011","10010011","10110011","00110011","00100011","11100011","00010011","00010011","10010011","11100011","00010011","10110011",
     "00110011","11100011","00010011","10010011","10010011","00010011","00010011","00010011","01101111","00010011","00010011","00010011","00010011","10010011","01100011","00000011",
     "00010011","00010011","10110011","10110011","10010011","00110011","11100011","00010011","00010011","00010011","10010011","00010011","10010011","11100011","00010011","10110011",
     "11100011","11101111","00010011","10010011","10010011","00000011","10010011","10010011","00110011","00100011","11100011","00010011","00110011","11100011","10000011","00000011",
     "00010011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","00010011","00010011","01100111","10010011","11101111",
     "10010011","00010011","11101111","10010011","00010011","11101111","10010011","00010011","11101111","01101111","00010011","00100011","00100011","00010011","00010011","10000011",
     "10000011","00000011","00000011","11101111","10010011","00000011","10000011","00010011","01101111","00010011","00100011","00100011","00100011","00010011","01100011","00010011",
     "10010011","10010011","10010011","00010011","01100011","01101111","00010011","00010011","10110011","10010011","11100011","10110011","00010011","10010011","10110011","01100011",
     "00110111","00010011","10010011","00010011","00010011","10110011","00010011","10010011","10010011","00110011","10010011","10010011","00110011","10010011","10010011","00010011",
     "00010011","00010011","00110011","00110011","00110011","00110011","00010011","00010011","10110011","00100011","10010011","00100011","11100011","00010011","10110011","11100011",
     "10110011","10010011","00000011","10010011","10010011","00100011","00100011","00100011","00100011","10000011","00000011","00010011","01100111","10010011","00010011","00010011",
     "10010011","01101111","00010011","01100011","10110011","10010011","10110011","10010011","00010011","00010011","00010011","10010011","10010011","00110011","10010011","01101111",
     "00010011","10010011","00010011","00010011","01100011","10000011","00010011","00010011","00110011","10110011","00010011","00110011","11100011","00010011","10010011","00010011",
     "10010011","00010011","11100011","00010011","10110011","11100011","01100111","00010011","01100111","01100011","00110011","00010011","10010011","00010011","00110011","10010011",
     "00010011","00110011","00010011","10010011","00000011","00010011","10010011","00110011","00100011","11100011","10010011","10110011","00110011","11100011","01100111","01100011",
     "10110011","10010011","00010011","10110011","00010011","00010011","10010011","10010011","00110011","10010011","00000011","10010011","00110011","00100011","11100011","10010011",
     "10110011","11100011","01100111","01100011","10010011","00010011","00110011","00110011","00100011","10010011","00010011","00010011","00000011","10000011","10010011","00010011",
     "00110011","00110011","00100011","11100011","10010011","00110011","11100011","01100111","01100011","00010011","00010011","00100011","00010011","00110011","00010011","10010011",
     "10110011","10010011","10010011","10010011","00100011","10010011","10010011","00010011","00000011","00000011","10010011","10110011","00110011","00110011","00100011","11100011",
     "10010011","10010011","11100011","10010011","00110011","00110011","10110011","11100011","00000011","00010011","01100111","01100111","01100011","00010011","00010011","00100011",
     "00010011","00110011","00010011","10010011","10110011","10010011","10010011","10010011","00100011","00010011","00010011","10010011","00000011","10000011","00010011","00110011",
     "10110011","00010011","10010011","00010011","10010011","10110011","10110011","00100011","11100011","10010011","10010011","11100011","10010011","00110011","00110011","10110011",
     "11100011","00000011","00010011","01100111","01100111","00010011","00010011","01100011","10010011","01100011","01100011","10010011","00010011","10110011","00100011","00100011",
     "00100011","00100011","00010011","11100011","01100011","01100111","10110011","10010011","10010111","10110011","01100111","00100011","10100011","00100011","10100011","00100011",
     "10100011","00100011","10100011","00100011","10100011","00100011","10100011","00100011","10100011","00100011","01100111","10010011","10010011","10110011","10010011","10110011",
     "01101111","10010011","10010111","10110011","10010011","11100111","10010011","10010011","00110011","00110011","11100011","01101111","00010011","00110111","00100011","00100011",
     "00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","00100011","10110111","00010011","00010011","10010011","00110011",
     "00010011","00100011","10110011","00010011","11101111","00010011","11101111","00100011","00010011","11101111","00100011","00010011","11101111","00100011","00010011","11101111",
     "00100011","00010011","11101111","01100011","00100011","00110111","00010011","10110111","00110011","10110011","00100011","10000011","01100011","00010011","01100011","10000011",
     "10000011","01100011","00000011","10110111","10010011","00100011","10010011","00100011","10000011","00110111","00010011","00110011","10110111","10110011","00010011","00010011",
     "10010011","00110011","00100011","00100011","00100011","10010011","00110011","01100011","00010011","00010011","00010011","00010011","00110011","00110111","00010011","00100011",
     "01100011","01100011","01100011","01100011","01100011","10010011","01100011","00110111","00010011","10110111","00110011","10110011","00000011","10000011","00000011","00100011",
     "11101111","10000011","01100011","10010011","00100011","10110111","10110111","10010011","10010011","10110011","10110011","00000011","00010011","10010011","10110011","10010011",
     "00100011","11101111","00000011","00100011","00100011","01100011","10010011","00010011","11101111","10000011","11101111","00100011","10010011","00010011","11101111","10000011",
     "11101111","00100011","01100011","00010011","11100011","11101111","11101111","11101111","11100011","10010011","10110011","00000011","10010011","10110011","00100011","00110111",
     "00010011","11101111","11101111","10110111","00110111","10010011","10110011","00010011","00110011","11101111","11101111","11101111","10010011","10110011","10110011","00010011",
     "00000011","10010011","10010011","00100011","11101111","10000011","10010011","00000011","11101111","10000011","10010011","00000011","11101111","10010011","00000011","11101111",
     "10110111","10010011","10010011","01100011","01100011","00110111","10010011","01100011","10110111","10010011","01100011","00110111","10110111","00010011","00010011","00110111",
     "11101111","00010011","00100011","00010011","10110111","10000011","10010011","10010011","01100011","10110111","10010011","10110111","10110011","10110011","00100011","00110111",
     "01101111","10000011","10110011","10010011","10110011","10110011","10000011","10110011","10010011","00010011","00000011","00010011","10010011","10010011","10010011","10010011",
     "01100011","00010011","10000011","10110011","10010011","10110011","10110011","10000011","00100011","10010011","01100011","00000011","01100011","10110111","10010011","10010011",
     "00010011","11101111","10000011","10010011","00100011","10000011","10110011","10010011","10110011","10110011","10000011","00010011","01100011","00000011","01100011","10000011",
     "10110111","10010011","00010011","11101111","00000011","10000011","00010011","00100011","10010011","11100011","10000011","00110011","00010011","00110011","00110011","00000011",
     "01100011","10000011","01101111","10000011","10000011","11100011","00000011","10010011","00100011","01101111","00110111","00010011","00110011","10110111","10110011","00000011",
     "10000011","00100011","11101111","10000011","00100011","00010011","11100011","00110111","00010011","00110011","10110111","10110011","00100011","00000011","10000011","00000011",
     "00000011","10000011","10010011","00110011","10010011","11101111","10000011","01101111","10110111","10010011","01100011","10110111","10010011","01100011","00110111","00010011",
     "00010011","00110111","00110111","11101111","00010011","00100011","00010011","01101111","10110111","10010011","10010011","00010011","11101111","10000011","10010011","10010011",
     "10010011","00100011","01101111","00110111","00010011","10110111","11101111","10000011","00110011","00110111","00010011","11101111","00110111","10010011","00010011","11101111",
     "10010011","00010011","11101111","10010011","00110111","00010011","11101111","00010011","00010011","10010011","00010011","11101111","01100011","00010011","10010011","11101111",
     "10010011","01100011","10000011","10000011","00110111","00010011","10110011","10010011","10010011","11101111","10110111","00110111","10010011","00010011","11101111","10110111",
     "00110111","10010011","00010011","11101111","10110111","00110111","10010011","00010011","11101111","00110111","10010011","00010011","11101111","10000011","10010011","01100011",
     "10000011","01100011","00110111","00010011","10110111","00110011","10110011","00010011","10110111","00100011","00110111","10010011","00000011","10110011","10010011","10110011",
     "10110011","00000011","10010011","00010011","11101111","00010011","10000011","00010011","00010011","11100011","10000011","10010011","01100011","10000011","01100011","00110111",
     "00010011","10110111","00110011","10110011","00010011","10110111","00100011","00110111","10010011","00000011","10110011","10010011","10110011","10110011","00000011","10010011",
     "00010011","11101111","00010011","10000011","00010011","00010011","11100011","10000011","10010011","01100011","10000011","01100011","00110111","00010011","10110111","00110011",
     "10110011","00010011","10110111","00100011","00110111","10010011","00000011","10110011","10010011","10110011","10110011","00000011","10010011","00010011","11101111","00010011",
     "10000011","00010011","00010011","11100011","00110111","10000011","00010011","00110111","00110011","00010011","00110111","00110011","10110111","01100011","10010011","10110011",
     "10010011","10110011","10110011","00000011","10010011","00010011","11101111","00010011","10000011","00010011","00010011","11100011","01100011","01100011","00110111","00010011",
     "11101111","00010011","11101111","00010011","10000011","00010011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011","00000011","10000011",
     "00000011","10000011","00010011","01100111","10010011","00100011","01101111","00110111","00010011","00110011","00110011","00010011","00100011","00100011","00010011","11100011",
     "01101111","00110011","10010011","00110011","00100011","11100011","01101111","00110011","00010011","10110111","00010011","00010011","00010011","00110011","00110111","00010011",
     "00110011","10110011","00100011","00100011","11100011","01101111","00110111","00010011","11101111","01101111","00100011","10010011","11100011","00010011","01101111","00110111",
     "00010011","11101111","01101111","00110111","00010011","11101111","00010011","01101111","10000011","10000011","10010011","00010011","10110011","11101111","10110011","00110111",
     "00010011","11101111","01101111","10010011","11100011","01101111","00110111","10110111","00010011","00010011","00110111","00110111","11101111","00010011","00100011","00010011",
     "01101111","00110111","10110111","00010011","00010011","00110111","00110111","11101111","00010011","00100011","00010011","01101111","00110111","00010011","11101111","00110111",
     "10010011","00110111","00010011","00100011","00010011","00010011","01101111","00010011","01101111","10010011","10010011","00010011","00010011","01100011","01100011","00110111",
     "01100011","10110111","01100011","10010011","10010011","00010111","00010011","00110011","00000011","10110011","00010011","00110011","01100011","00110011","10110011","10110011",
     "00110011","00110011","00010011","00110011","10010011","10010011","10010011","00110011","10110011","00010011","00110011","01100011","00110011","10010011","01100011","01100011",
     "00010011","00110011","00110011","00010011","00010011","00110011","10110011","00010011","00110011","01100011","00110011","10010011","01100011","00010011","01100011","00010011",
     "00010011","00110011","10010011","01100111","01100011","00010011","10110011","00110111","01100011","10110111","01100011","10010011","10010011","00010111","00010011","00110011",
     "10000011","10110011","10010011","10110011","01100011","10010011","00110011","00010011","10010011","10010011","10010011","00110011","00110011","10110011","00010011","10110011",
     "01100011","10110011","00010011","01100011","01100011","00010011","10110011","00110011","00010011","00010011","10110011","10110011","10010011","10110011","01100011","10110011",
     "10010011","01100011","00010011","01100011","00010011","00010011","00110011","01100111","01100011","10110111","01100011","10110111","01100011","00010011","00010011","10010111",
     "10010011","10110011","00000011","00010011","00110011","00110011","01100011","01100011","00110011","00010011","10010011","01100111","10010011","00010011","01100111","10010011",
     "01100011","00010011","00010011","01101111","00010011","10010011","11100011","10010011","10010011","01101111","00010011","10010011","11100011","10010011","10010011","01101111",
     "10110011","00110011","00010011","00110011","00110011","10110011","00110011","10010011","10010011","00110011","10010011","10110011","10110011","10010011","10110011","01100011",
     "10110011","00010011","01100011","01100011","00010011","10110011","10110011","00110011","10010011","10010011","10110011","00110011","00010011","00110011","01100011","00110011",
     "10010011","01100011","01100011","00010011","00110011","10010011","00110011","10110011","01101111","10110011","10110011","10110011","00110011","00010011","10110011","10010011",
     "10010011","00110011","00110011","00110011","10010011","00110011","00110011","10110011","00010011","10110011","01100011","10110011","00010011","01100011","01100011","10010011",
     "10110011","10110011","00110011","00010011","00010011","10110011","00110011","10010011","10110011","01100011","10110011","00010011","01100011","01100011","00010011","10110011",
     "10010011","00110111","10110011","00010011","10110011","10010011","00110011","00010011","10110011","10110011","10110011","00010011","00110011","10110011","10110011","00110011",
     "01100011","00110011","10010011","00110011","01100011","01100011","00010011","10010011","01100111","00110111","00010011","10110011","10010011","10110011","00110011","10110011",
     "11100011","00010011","10010011","01100111","00010011","00010011","01101111","10010011","10010011","01101111","10010011","10010011","01101111","10010011","00010011","01100111",
     "00010011","00010011","01101111","00010011","01101111","00010011","01101111","10010011","01101111","00010011","01101111","00010011","00110011","01101111","00010011","10110011",
     "01101111","10110011","10010011","10110011","01100011","10010011","01100011","10010011","00010011","01100011","00010011","10010011","01100011","01100011","10010011","10010011",
     "00000011","10010011","10010011","00100011","11100011","10010011","10110011","10010011","10010011","00110011","10110011","01100011","01100111","00010011","11100011","10000011",
     "00010011","10010011","10100011","11100011","01100111","10000011","00010011","10010011","10100011","10010011","11100011","10000011","00010011","10010011","10100011","10010011",
     "11100011","01101111","10000011","10000011","10000011","00000011","10000011","00000011","00000011","00000011","10010011","00100011","10000011","00100011","00100011","00100011",
     "00100011","00100011","00100011","00100011","00010011","00100011","11100011","01101111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
  signal ram_symbol1 : ram_type := (
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00101110","00101100","00101010","00101000","00100110","00100100","00100010","00100000",
     "00101110","00101100","00101010","00101000","00100110","00100100","00100010","00100000","00000001","01000000","00100000","00100010","00100011","00100011","00100101","00100101",
     "00100110","00100110","00100111","00100111","00101000","00101000","00101110","00101110","00101111","00101111","00000001","00000000","00100001","10000001","00010001","00000001",
     "00100101","00000101","10000101","00001000","00100000","00000101","11110000","01110101","00000101","00000001","01110101","10000101","00001110","00100110","00000101","00100000",
     "10000000","00100101","11110000","00000001","00010101","00000101","00010000","00100101","00000101","00010000","01010000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00011111","00011110","00011110","00011111","00011111","00011110","00101111","00101111","00101111","00101111","00101111","00101111","00101111","00101111","00101111","00101111",
     "00101111","00101111","00101111","00101111","00101111","00101111","00101111","00110110","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010",
     "00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110000","00110010",
     "00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110100","00110010","00110001","00110110","00110010","00110010","00110010","00110010","00110110",
     "00110010","00110010","00110010","00110010","00110010","00110001","00110001","00110010","00110010","00110000","00110010","00110000","00110010","00110010","00110100","00110010",
     "00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010",
     "00110010","00110010","00110010","00110010","00110010","00110010","00110000","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110100",
     "00110010","00110001","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110010","00110001","00110001","00110010",
     "00110010","00110000","00110010","00110000","00110010","00110010","00110000","00110001","00110101","00111001","01100100","01101000","01101100","01110000","01110100","01111000",
     "00000000","00110001","00110101","00111001","01000100","01001000","01001100","01010000","01010100","01011000","00000000","01001110","00111110","01100101","01110011","00100000",
     "01100011","01101111","01110101","01101110","01110100","00100000","00000000","01100101","01110011","00100000","01100011","01101110","01101111","01100001","00101000","01101001",
     "01100001","01101110","00100000","01110011","01111001","01101011","01101111","01110100","00101110","00001010","01001110","01010110","00100000","00100000","01101111","01100100",
     "01101101","01110011","01101100","01101000","01110100","01101001","01100111","01110000","00101110","00000000","01110100","00100000","01100101","00000000","01101011","01110010",
     "01101101","01100101","01101110","01110010","01110100","00100000","00100000","01100101","01101011","00000000","01101011","01101100","01110100","00100000","00100000","01100001",
     "01100101","01100110","01100011","01101101","00101110","01110010","01101100","01100101","01100001","01101110","01101110","01110010","01110100","00100000","00100000","01100101",
     "01101011","00000000","01001011","01110010","01101101","01100101","01101110","01110010","01110100","00100000","00100000","01100101","01101011","00000000","01001011","01101100",
     "01110100","00100000","00100000","01100001","01100101","01100110","01100011","01101101","00101110","00100101","01010010","00100001","01110011","01110010","01111000","01111000",
     "01110011","01101100","01100101","00100101","00001010","00100101","01010010","00100001","01110100","00100000","00100000","00110000","00101101","01101111","00100000","00110000",
     "00110100","00000000","00100101","01010010","00100001","01100001","01100011","00110000","00110100","00100000","01110101","01100010","01111000","01111000","01101111","01100001",
     "01010011","00100000","00111010","01110101","01101111","00100000","01101011","00100000","00111010","01110101","01101111","00100000","01100101","01100101","00111010","00001010",
     "01110100","01110100","01110011","01100011","00111010","00001010","01010010","00100001","01110011","01111000","01110100","01101111","01110100","01100001","00110001","01100101",
     "01100110","01100001","01101100","01110010","01101100","00000000","01110100","01110100","01110011","00100000","00111010","01110101","01000011","00110011","00000000","01101111",
     "01101100","01110110","01101001","00111010","00001010","00111110","01100110","01110100","01100101","01100001","01101001","00000000","01101111","01101100","01100110","01110011",
     "00111010","00001010","01010100","00000000","01100101","01111001","01100011","01101111","00111010","00001010","01100101","01110010","00100000","00100000","00111010","00100101",
     "00001010","00100101","01110010","01110011","00100000","00100000","01111000","01111000","00100101","01110010","01110100","00100000","00100000","01111000","01111000","00100101",
     "01110010","01100001","00100000","00100000","01111000","01111000","00100101","01110010","01101110","00100000","00100000","01111000","01111000","01101111","01100011","01110000",
     "01110100","00100000","01101001","01100101","01010011","01010010","01001101","01100100","01110010","01101110","01100100","01110000","01101001","01110010","01110011","00000000",
     "01110010","01110011","01110100","01100101","00000000","01100001","01110100","01101100","01110100","01110000","01110100","00100000","00100000","01110011","01100101","01110110",
     "01100101","01110000","01110011","01101111","01110010","01101001","01110010","01101100","01101111","00100000","01110111","01101100","01101111","00001010","01110100","01100011",
     "01100101","00000000","01110100","00000000","01001011","01001011","01001011","01001011","01001100","00011101","00011101","00011101","00011101","00011101","00011101","00011101",
     "00011101","00011101","00011101","00011101","00011101","00011100","00011100","00011100","00011101","00110000","00101101","00000000","01010100","00101011","00000000","01010100",
     "01100101","00000000","00110100","00101101","00000000","00101110","01100101","00000000","00101110","01100101","00000000","00111000","00111000","00000000","00110000","00101101",
     "00000000","00110101","00110100","00000000","00110001","00110101","00000000","00110001","00110111","00000000","00110000","00110100","00000000","00110000","00000000","00110010",
     "00000000","00111000","00000000","00110001","00000000","00000001","00000011","00000100","00000100","00000101","00000101","00000101","00000101","00000110","00000110","00000110",
     "00000110","00000110","00000110","00000110","00000110","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",
     "00000111","00000111","00000111","00000111","00000111","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000111","11100110","00010111","10000111","00010101","00000101","00100111","10000000","00100111","10100101","10000000","10100101","10000000","10100101",
     "10000000","00100111","10100101","10000000","10100101","10000000","00000101","10000000","01000110","11110110","01010111","11010111","10001100","10100110","10000110","11000111",
     "10010111","11010111","11000111","01110111","01010110","11010111","00001100","10100111","00000111","11000111","10010111","11010111","11000110","11110110","01010111","11010111",
     "10001100","10100110","10000110","11000111","10010111","11010111","11000111","01110111","01010110","11010111","00001100","10100111","00000111","11000111","10010111","11010111",
     "11000110","11110110","01010111","11010111","10001100","10100110","10000110","11000111","10010111","11010111","11000111","01110111","01010110","11010111","00001100","10100111",
     "00000111","11000111","10010111","11010111","11000110","11110110","01010111","11010111","10001100","10100110","10000110","11000111","10010111","11010111","11110110","11010101",
     "10001100","10100111","10000111","01000111","10010101","01010101","10000000","11000110","01110110","01110110","11010111","11010111","00001100","10100110","00000110","11000111",
     "10010111","11010111","11000111","01110110","11010111","11010111","00001100","10100110","00000110","11000111","10010111","11010111","11000111","01110111","11010110","11010111",
     "00001100","10100111","00000111","11000111","10010111","11010111","11000110","01110110","11010111","11010111","00001100","10100110","00000110","11000111","10010111","11010111",
     "11000111","01110111","11010110","11010111","00001100","10100111","00000111","11000111","10010111","11010111","11000110","01110110","11010111","11010111","00001100","10100110",
     "00000110","11000111","10010111","11010111","11000111","01110111","11010110","11010111","00001100","10100111","00000111","11000111","10010111","11010111","11110111","11010111",
     "00001100","10100111","00000111","11000111","10010111","11010111","01010101","11000110","01110111","01110110","01010110","11010101","00001100","10100111","10000111","01000101",
     "00010101","01010101","11000110","11110110","01010111","01010101","10001100","10100110","10000110","01000101","00010101","01010101","01000111","11110111","01010110","01010101",
     "10001100","10100111","10000111","01000101","00010101","01010101","01000110","11110110","01010111","01010101","10001100","10100110","10000110","01000101","00010101","01010101",
     "01000111","11110111","01010110","01010101","10001100","10100111","10000111","01000101","00010101","01010101","01000110","11110110","01010111","01010101","10001100","10100110",
     "10000110","01000101","00010101","01010101","01000111","11110111","01010111","01010101","10001100","10100111","10000111","01000101","00010101","01010101","01110111","01010101",
     "10001100","10100111","10000111","01000101","00010101","01010101","10000000","11001000","01110110","00010111","01111000","01010111","11010110","11010111","00001100","10100101",
     "10000101","11000111","10010111","11010111","11000110","01110101","11010111","11010110","10001100","10100101","10000101","11000111","10010111","11010111","11000110","01110110",
     "11010101","11010111","00001100","10100110","00000110","11000111","10010111","11010111","11000101","11110101","11010110","11010111","10001100","10100101","10000101","11000111",
     "10010111","11010111","11000110","01110110","11010101","11010111","00001100","10100110","00000110","11000111","10010111","11010111","11000101","11110101","11010110","11010111",
     "10001100","10100101","10000101","11000111","10010111","11010111","11000110","01110110","11010110","11010111","00001100","10100110","00000110","11000111","10010111","11010111",
     "11110110","11010111","00001100","10100110","10000110","11000111","10010111","11010111","01010111","11000110","11110110","01110111","01010110","11010111","10001100","10100110",
     "10000110","11000111","10010111","11010111","11000110","01110110","01010110","11010111","00001100","10100110","00000110","11000111","10010111","11010111","11000110","11110110",
     "01010110","11010111","10001100","10100110","10000110","11000111","10010111","11010111","11000110","01110110","01010110","11010111","00001100","10100110","00000110","11000111",
     "10010111","11010111","11000110","11110110","01010110","11010111","10001100","10100110","10000110","11000111","10010111","11010111","11000110","01110110","01010110","11010111",
     "00001100","10100110","00000110","11000111","10010111","11010111","11000110","11110110","01010111","11010111","10001100","10100110","10000110","11000111","10010111","11010111",
     "11110110","11010111","10001100","10100111","00000111","11000111","10010111","11010111","01010101","11000101","01110111","00010110","11110101","11010110","01010110","11010101",
     "10001100","10100111","10000111","01000101","00010101","01010101","01000110","01110110","01010111","01010101","00001100","10100110","00000110","01000101","00010101","01010101",
     "01000111","11110111","01010110","01010101","10001100","10100111","10000111","01000101","00010101","01010101","01000110","01110110","01010111","01010101","00001100","10100110",
     "00000110","01000101","00010101","01010101","01000111","11110111","01010110","01010101","10001100","10100111","10000111","01000101","00010101","01010101","01000110","01110110",
     "01010111","01010101","00001100","10100110","00000110","01000101","00010101","01010101","01000111","11110111","01010111","01010101","10001100","10100111","10000111","01000101",
     "00010101","01010101","01110111","01010101","10001100","10100111","10000111","01000101","00010101","01010101","11010111","01000111","01110111","11110111","11010110","01010101",
     "00001100","10100111","00000111","01000101","00010101","01010101","01000110","11110110","11010111","01010101","10001100","10100110","10000110","01000101","00010101","01010101",
     "01000111","01110111","11010110","01010101","00001100","10100111","00000111","01000101","00010101","01010101","11000110","11110110","11010111","01010101","10001100","10100110",
     "10000110","01000101","00010101","01010101","01000111","01110111","11010110","01010101","00001100","10100111","00000111","01000101","00010101","01010101","11000110","11110110",
     "11010111","01010101","10001100","10100110","10000110","01000101","00010101","01010101","01000111","01110111","11010111","01010101","00001100","10100111","00000111","01000101",
     "00010101","01010101","01110111","01010101","00001100","10100111","10000111","01000101","00010101","01010101","10000000","11000110","01110111","00010111","01110110","11010111",
     "01010110","11010101","00001100","10100101","10000101","01000101","00010101","01010101","01000110","11110110","01010101","01010110","00001100","10100101","10000101","01000101",
     "00010101","01010101","01000110","11110110","01010110","01010101","10001100","10100110","10000110","01000101","00010101","01010101","01000110","01110110","01010110","01010101",
     "00001100","10100110","00000110","01000101","00010101","01010101","01000110","11110110","01010110","01010101","10001100","10100110","10000110","01000101","00010101","01010101",
     "01000110","01110110","01010110","01010101","00001100","10100110","00000110","01000101","00010101","01010101","01000110","11110110","01010111","01010101","10001100","10100110",
     "10000110","01000101","00010101","01010101","01110110","01010101","10001100","10100111","00000111","01000101","00010101","01010101","11010111","01000111","01110111","11110111",
     "11010110","01010101","00001100","10100111","00000111","01000101","00010101","01010101","11000110","11110110","11010111","01010101","10001100","10100110","10000110","01000101",
     "00010101","01010101","01000111","01110111","11010110","01010101","00001100","10100111","00000111","01000101","00010101","01010101","01000110","11110110","11010111","01010101",
     "10001100","10100110","10000110","01000101","00010101","01010101","01000111","01110111","11010110","01010101","00001100","10100111","00000111","01000101","00010101","01010101",
     "01000110","11110110","11010111","01010101","10001100","10100110","10000110","01000101","00010101","01010101","01000111","01110111","11010111","01010101","00001100","10100111",
     "00000111","01000101","00010101","01010101","01110111","01010101","00001100","10100111","10000111","01000101","00010101","01010101","10000000","00000101","10000000","00000001",
     "00101010","00100100","00101110","00101100","00101000","00100110","00100010","00100000","00101110","00101100","00101010","00101000","00100110","11111000","00000100","00001010",
     "00000110","00011000","10001000","11111101","00010000","11110110","11111110","00001100","00001100","11110110","11111101","00000110","11001000","11110110","00011010","11110111",
     "00000011","10000110","10000110","00000011","10001100","00000111","00001100","00000111","10110111","10000110","10010100","00000111","00001110","00001001","00001100","00001001",
     "00000100","10001010","11010100","00001010","10001011","00001011","00010110","01011100","00000110","10000101","00000101","00100110","00100000","00100011","10000100","00001011",
     "00001011","00000110","10000000","10000100","10001010","00000111","00000000","00000111","00001100","00011100","01010000","11001010","01011010","11111010","00001101","10001011",
     "10000101","00000110","00000101","00001011","00100000","10000100","00001011","11011110","10001010","10000101","10000110","00000101","00100000","10000100","00000110","10000111",
     "00000101","00000111","01000101","00000111","10000111","00001111","10000111","00000110","01000010","10000100","01010100","11000111","11010111","11110100","00000100","10000101",
     "00000110","00000101","00100000","10000100","00100000","00100100","10000101","00101001","00100100","00101001","00101010","00101010","00101011","00101011","00101100","00101100",
     "00101101","00101101","00000001","10000000","11110111","00001110","11110110","00001100","11111101","00001010","11110000","00011000","10001000","11110000","00000011","11110000",
     "00000101","10000110","00000011","10010100","00001001","00000100","00000000","10001001","11110111","00001001","00001000","10000101","10001100","10000111","11000111","11010101",
     "00001111","01111100","11110000","10000110","00000011","11110000","00000111","10000000","00000111","10000000","10000100","11110000","10000110","11110000","00000111","10000000",
     "10000100","11110000","10001011","10001011","11110000","00000111","10001011","10001011","11110000","00000111","00000000","00000111","00100111","11010111","11110111","10001010",
     "00100000","10000000","00000111","00100111","11010111","11110111","10001010","00000111","00100000","11110000","00000001","00100100","00100110","00100100","00100010","00100000",
     "00101110","00101100","00101010","00101000","00100110","00100010","00100000","00101110","00101010","00101100","00101110","00100000","00100010","00100100","00100110","01000111",
     "00001100","00101010","10000000","00001001","00011011","00011010","00011001","00000100","00001011","10001011","00001010","10001001","00011010","00000111","10001010","00000000",
     "01000111","00001011","00000100","10010100","00000000","01000110","10000010","00000110","00000101","00000111","00001000","00000110","10000010","00100111","11010111","11110111",
     "10001010","00000101","00100000","00001001","01000110","10011110","00100000","00100100","00100100","00101001","00101001","00101010","00101010","00101011","00101011","00101100",
     "00101100","00101101","00101101","00000001","10000000","00100111","11010111","11110111","10001010","00100000","11110000","01000101","00000110","00000111","10000111","01110111",
     "00000100","11101000","00010111","00000111","00100111","00000000","11100111","10000100","01000101","00000100","10000111","01110111","11111100","10000111","01110111","00000110",
     "11111010","00000111","00000110","10001110","00000110","00000111","10001000","11110110","00000101","00001010","10000110","01110110","00000101","01101100","00010110","00000110",
     "00100110","00000000","11100111","10000100","11110000","11100111","10000100","11110000","11100111","10000100","11110000","11100111","10000100","11110000","11001000","00000101",
     "10001100","00000110","01110110","01100100","00010101","00010110","00000101","00000110","00100110","00000000","11000101","00000110","10000101","10000111","01110111","01110100",
     "00000111","10001100","00000100","00000111","11110000","00000110","00000110","10010111","00000110","10000100","10010110","10000110","11000101","10000110","10000111","01110111",
     "01111110","11110000","00100110","00000100","01000101","00001100","11011100","00000110","11100111","11110000","10001100","11100111","00000110","00000101","00100101","00001100",
     "00000101","11110000","11000111","00001011","10000100","10010000","11110000","10001100","00000110","11110000","10001100","00100100","00001100","00000000","01000110","00001000",
     "00000110","00000110","00000000","00000101","10001000","00000110","01000101","10011000","11110111","00000100","10001010","01010010","00000111","00000110","00110111","00110110",
     "10000111","01000111","01000110","10110111","01100111","11000111","11110111","10000110","01100111","11110111","10010000","11110101","00000111","00000111","10000101","10100110",
     "00000111","10000111","00101110","10011000","11110111","00000100","00000110","00000111","10000110","01000101","10000101","00000000","11011110","01000101","10000111","00000000",
     "11010110","01000111","00000001","00001011","10000100","11011110","10000100","00000101","10000110","00000101","00100000","00001011","11000111","10010000","11110000","10001100",
     "00000110","10000010","00100101","00000110","00001100","11110000","10001100","00000110","11110000","10001100","11110111","10000100","10000010","00100111","00000111","00001100",
     "00000000","10000100","01010100","10000110","00000101","00000101","00100000","11000111","00001011","10011000","11110000","10001000","10001100","00000111","00000111","00001010",
     "00000000","11001000","00011110","00001011","00000000","01000110","10010010","00000101","11110000","00000111","00001000","00010110","00000111","00000101","00010111","00000111",
     "01000101","00000111","10000110","01110110","01111110","00000100","11110000","00100111","11000101","00001100","01000110","01010110","01110111","10000100","11110000","00001000",
     "11100111","00000101","00000110","10000110","00000000","00000110","00100111","11100111","00001100","10011000","00010110","00000110","01001000","01000101","01001110","01000011",
     "01001000","01000101","01010011","01010010","01011111","01011111","11011110","01111000","01110101","01111110","01110011","11111000","11010111","00001000","00000101","00000011",
     "00000010","00001111","00001110","00001111","00000011","00001110","00001000","01000100","01001100","11000011","11000010","11001111","01001110","01001111","01000011","11001110",
     "11001000","00000101","01000101","00000111","11110101","00001100","00001101","00001110","00000000","00000001","00000011","00001100","00001101","00001110","00001111","00001111",
     "00000000","00000001","00000010","00000010","00000111","00000011","01000111","11110111","10000100","00000100","10011010","00000111","11010000","10000100","00000110","00000101",
     "00000101","00100110","00100000","00000110","00000101","00000101","00110000","00100110","00000111","11000111","10000100","00001011","10010010","11110000","00000110","00100111",
     "00001100","10011000","10000110","11110000","10001100","00000110","11110000","00100111","00001100","01000110","00000100","00000101","11011110","00000101","01101000","00001000",
     "00000101","00000100","00000011","01000110","11000101","10000110","01000110","00001100","10000110","01000101","11100110","00001100","10000110","01000110","00000101","00000011",
     "00000100","00000101","01000110","00000101","00001000","00000100","00000000","00001000","01010110","00001000","00001000","00001110","00001110","00000101","01100011","01000110",
     "01001000","10000110","01000110","00000100","10000110","01001000","01100110","00000101","10000110","01000101","00000110","00000110","10000100","00000100","00000101","01000110",
     "10000101","00000101","00000100","00000101","00001100","00001000","01010010","00001000","00001000","00001110","00001110","00000101","01100011","01000110","01001000","10000110",
     "01000110","00000100","10000110","01001000","01100110","00000101","10000110","01000101","00000110","00000110","10000100","00000100","01000111","00000110","00000101","00000110",
     "10000100","00000110","00001000","00000101","01010110","00000101","00001000","00000011","00000011","00000110","01101000","01000111","11000101","10000111","01000111","00000100",
     "10000111","01000101","11100111","10000101","10000111","01000101","00000111","00000111","00000100","00000100","11110111","10001100","10011010","01011000","10001101","00000101",
     "00000110","00000101","00100110","00100000","00100110","00001011","00000110","10000110","10001100","00000101","00000110","00000101","00100110","00110000","00100110","00000111",
     "00001011","01010010","00000110","00000110","00001011","10000111","10000111","00001111","00000111","01000110","11000111","10000100","10010010","11110000","11100111","00000101",
     "10001100","00100101","00000110","00001100","11110000","00100111","11100111","00001100","11110000","00000111","00001011","10000111","00000000","11000111","10000100","00001011",
     "10011010","11110000","11100111","00000110","11110000","01010100","10000110","00000101","00000101","00001011","00100000","00000100","11110000","10000100","11110000","10001101",
     "11010000","10001101","00000101","10000110","00000101","00100110","00100000","00100110","00001011","10000110","10000110","11110000","00000110","00001100","00000100","00000101",
     "01000110","00000101","00001000","00000100","00000101","00010100","00000110","00000110","00000101","00000100","00000100","00000101","01000110","10000101","00000101","00000100",
     "00000101","00011000","00000110","00000110","00000101","00000100","00000100","00000110","01000111","00000101","00000110","10000100","00000110","00011100","00000111","00000111",
     "00000110","00000100","00000100","11110000","10000111","00000110","10000100","00000110","00000101","00000101","00100110","00110000","00100110","00001100","00000111","11010100",
     "00000101","00000110","00000110","00000111","00000111","00000111","00001111","10000111","11000110","11110000","00001001","00001011","11110000","10000100","11110000","00000101",
     "01011100","00001000","01000101","00001000","10001000","00000101","10000101","01000101","01100110","10000100","11110000","00000101","01011000","00001000","01000101","00001000",
     "10001000","00000101","10000101","01000101","01100110","10000100","11110000","00000101","11011000","00000101","01000101","00001000","00001000","00000110","10000101","11000101",
     "01100111","00000100","11110000","00000101","11010110","00001000","01000101","00000101","00000100","00000011","10000101","01000101","01100110","00001100","11110000","00000101",
     "00000100","00000011","11110000","11110100","10000110","00000100","11110000","00100111","00000111","00001100","00000000","10000100","11000111","00001011","10011110","11110000",
     "00000110","11110000","00000111","00000100","01000111","00001011","00001111","00011000","11110000","10000111","10000110","10001100","11110000","00000001","00101000","00101110",
     "00101100","00101010","00100110","00010100","01010111","11110111","01111001","10011110","10000100","01010101","11110101","10010111","01110111","11100101","00001001","11010111",
     "00001100","00000110","00001010","00010101","01010101","00001001","10000101","01111001","01110100","11100000","01100100","10011100","01100100","10010000","00100000","00100100",
     "00000101","00100100","00101001","00101001","00000001","10000000","00000110","10000111","11010100","00000111","10010110","10010110","10100101","10100101","01110111","00010000",
     "11010111","00011001","01011001","10010100","10011111","11010111","11110000","10000110","10000101","00010000","11010111","00011001","01011001","10010000","11010111","10011110",
     "11110000","00000001","00101010","00101000","00100100","00101110","00101100","00100110","00010100","10001001","00000100","01010111","11110111","01111010","10011100","01010101",
     "11110101","10010111","01110111","11100101","00001001","01010111","00000000","00000110","00000000","00010101","01010101","00001010","10000101","01111010","01110100","11100000",
     "01100100","10011100","01100100","10010000","00010100","01010111","11110111","01111001","10011010","01010101","11110101","10010111","01110111","11100101","11010111","00000000",
     "00000110","00000010","00010101","01010101","00001001","10000101","11111001","01110100","11100000","11100100","10011100","01100100","00010000","00100000","00100100","00000101",
     "00100100","00101001","00101001","00101010","00000001","10000000","00000110","10000111","11010100","00000111","10010110","10010110","10100101","10100101","01110111","00010000",
     "11010111","00011010","01011010","10010100","10011111","11010111","11110000","00000110","10000111","11010100","00000111","10010110","10010110","10100101","10100101","01110111",
     "00010000","11010111","00011001","11011001","10010100","10011111","11010111","11110000","10000110","10000101","00010000","11010111","00011010","01011010","10011110","11010111",
     "10011110","11110000","10000110","10000101","00010000","11010111","00011001","11011001","10011100","11010111","10011110","11110000","00001010","00010101","10010111","00000101",
     "10000000","00010111","10010111","01010111","01010111","11110111","11100111","00010000","10010111","10010111","01010111","01010111","11110111","11100111","10010000","00010101",
     "10010111","00000101","10000000","10010111","00010000","10010111","00010001","10000000","00000001","00101100","00101110","00101100","00101010","00101000","00100110","00100100",
     "00100010","00100000","00101110","00101010","00101000","00100110","00011000","00101010","00001100","00100100","01011000","00100110","00000110","00001110","00000101","00001000",
     "00100111","01110110","00101010","11001000","00001110","00100111","10000110","00000111","00010111","00011100","00000000","10100111","00100110","00010111","00000110","10100111",
     "10010110","00000110","00000000","00000110","00000100","00100111","00100000","00011000","10001000","10100111","00000101","00010101","00010111","01010101","01110110","10001100",
     "01010111","01110111","00000111","00011000","01011000","10100110","10001100","10100111","10100000","00100111","10100000","00100000","00100111","11001010","10001011","00010111",
     "11010111","00100110","00000110","00010110","01010110","10010110","00010111","10000111","00000111","10010111","11010111","00101110","01001100","00100111","00000100","10101001",
     "10100111","00100110","10100010","00100010","10100111","00100111","10100000","00100111","00100000","11001110","10100111","00100111","10010111","10001010","10100100","10010110",
     "00100100","10000010","00100111","00100101","10010101","11100000","10100100","00101110","10010100","00100100","10100111","00100111","00000011","00100010","10100111","10100010",
     "00001000","00100000","10100000","00001110","00000100","00001111","00001110","00000110","00000111","10100110","10000111","10000110","00011010","00000111","00000111","00000110",
     "10000100","10001100","00001110","00001100","00100101","00100101","10010110","10011000","01011000","01011000","11110110","11100110","10010000","00010110","00011110","10011000",
     "01011000","11110110","01011000","11100110","00010000","10010110","10000110","01010100","00000110","00100100","00000110","10000100","10100000","10001000","10011000","00001100",
     "00001100","00000110","00000110","00100100","10010000","10000100","10001000","11110000","10100111","00100111","11000111","10001110","10100100","10010110","00100100","10010110",
     "11110000","00000110","10000111","00100111","11110000","00010010","10100000","00001110","00010011","10000000","10000100","00001110","00001000","00000100","11110000","00001000",
     "00100111","00000111","01000111","10011100","11110000","10100111","00100110","01000111","00000010","10100111","10010110","11110000","10100111","00000111","10011110","00000111",
     "01011110","01110111","00000111","00011000","01011000","11110000","10100100","00000100","10100111","00100101","10010101","11100000","00100100","00101110","00010100","00100000",
     "00100100","00100100","00101001","00101001","00101010","00101010","00101011","00101011","00101100","00101100","00101101","00101101","00000001","10000000","00100110","00101110",
     "01011010","00000000","00000111","00100100","00000111","00101100","00001101","00001001","00000100","00101000","00001010","00100111","00001101","00001011","10000111","00101000",
     "10101101","10001011","10000110","00100111","10011000","00101100","10001000","10001000","10000110","00101010","10101001","10010100","11110111","11111011","10011000","11010101",
     "11110101","10010111","11110111","11100101","01010111","00000110","00000000","10010101","01010101","10001011","10000101","11010000","01111011","11111000","01101000","00011100",
     "11101000","10010000","10011010","11110111","11110100","10011000","11010101","11110101","10010111","11110111","11100101","01010111","00000010","00001100","10010101","01010101",
     "10000100","10000101","11010000","11110100","11111000","11101000","00011100","11101000","10010000","00000100","01010010","10000111","10101101","10001100","00000100","00100000",
     "10001001","10011100","10001010","10001100","10000111","10001100","10101101","00010000","10000100","10001001","11110000","00000111","10001011","00101101","11110000","10001101",
     "10010110","00100111","00100000","00000111","00000010","00100111","10010111","00100100","00011100","00100000","00000000","00100101","10000110","00010000","01010111","00010100",
     "11010100","10010110","01010111","00011110","11110000","00000110","10000111","11010100","00000111","00010110","00010110","00100101","00100101","01110111","00000000","01010111",
     "00010100","11010100","10010100","00011111","01010111","11110000","00100101","10000110","00010000","01010111","00011011","01011011","10010110","01010111","00011110","11110000",
     "00000110","10000111","11010100","00000111","00010110","00010110","00100101","00100101","01110111","00000000","01010111","00011011","01011011","10010100","00011111","01010111",
     "11110000","00100101","11110000","00100111","00000000","00000111","01010101","10100000","10000111","10001000","10000110","10001000","00000101","00011111","10001111","10100010",
     "00010001","10100111","00011111","00001111","00010000","00000011","11110010","00001000","10100111","01110100","10100100","10100000","10100110","00000111","11000111","00010010",
     "00010011","10100111","00001010","00010011","10000010","11010011","00001000","11000010","10001110","01111000","00001110","11110100","10010011","01010011","01000111","10010111",
     "11110111","01110011","10100000","11100111","10100000","10010111","10100010","01100111","00010000","00010001","10100111","10001000","00000110","10001000","00010100","00100111",
     "10001010","00000111","01010101","01000011","00000110","00000011","00101000","11110000","10010001","00100111","10000110","00100111","10010100","00001111","00000011","10000111",
     "00001000","00000101","00001111","00001111","10000101","00000111","00100101","00000111","00000100","00011010","10000110","10000110","00000111","00001100","00001100","10001010",
     "10100011","10101110","00011000","00010101","01010101","01010101","01111000","01101000","00010000","00011000","00010010","00011110","11011110","01111000","11011110","01101000",
     "00010000","00010101","00000101","01010010","10001000","10100111","00000110","10000100","10100000","00001000","00011000","00001010","10001010","10001000","00000110","10100111",
     "10010000","00000101","00001000","11110000","10001000","00000111","10100110","11110000","10010110","10100000","00000110","10011111","10010110","00100000","00000000","10011000",
     "01011000","00000111","10010111","11110111","01001000","11100111","11110111","10010001","00100111","10000110","00100111","10010110","11110000","10000101","10000000","10100111",
     "00001000","10000110","11110000","00001000","10000110","11110000","00101000","00001000","11110110","10100111","00000111","01110000","00100000","00100111","00100000","00100000",
     "10100111","00000101","00100010","10000111","10100000","10010111","00100111","10010000","10010111","10010001","10000000","00001000","00000101","10000000","00100111","00100110",
     "00000111","00100110","00000101","10100010","00100010","10100110","10100110","10100000","00100000","10000000","10100111","00100110","00100010","10100111","10100010","00100000",
     "10100000","10000000","10010111","01001000","00000100","00100111","10010111","10011010","00000000","00100111","10010111","10000110","00100101","00011000","10000000","00001110",
     "00100111","10010111","11000111","10011010","00000000","00100111","11000111","10001000","00100101","00011000","11110000","10000000","10000000","10000000","00000000","00000111",
     "00000000","10000101","00100111","00100000","00000111","10011000","10000000","00000100","00000001","00101010","00101000","00100110","00100100","00100000","00100110","00100100",
     "00100010","00100000","00101110","00101100","00100010","00001011","10001011","00001100","00001010","00001101","00001010","00001100","00001001","00001011","10001100","00000100",
     "00000100","00100100","10000100","00000100","10011010","10001001","10001110","10001110","00001100","00100101","00100101","00000110","10000000","01010010","00000111","00100100",
     "10001001","00000100","00100000","10001001","10010110","10001010","00001100","00000111","10001001","00100100","00010000","10001011","10001001","11110000","00000111","10000100",
     "00101010","11110000","00001010","00010110","00100000","10001010","10011010","00010110","00100000","00000000","00100000","00100100","00000101","00100100","00101001","00101001",
     "00101010","00101010","00101011","00101011","00101100","00101100","00101101","00000001","10000000","00100000","00000000","00000101","00000101","10000000","00100111","00000110",
     "00000110","00101010","00101000","00000111","10100000","01000110","10100100","00000111","10000110","10100000","00000110","10100010","00000111","10100000","10000000","00000111",
     "10100111","00100111","10100110","10100100","10000000","00100111","00100111","10100101","00100101","10100111","00100111","10000101","10110101","10000111","10000101","10000000",
     "00000001","00000110","00000110","00100110","00010000","00100000","00000001","10000000","00000001","00100100","00000100","00010101","00000101","00000101","00100110","11100000",
     "00010101","00000101","00000101","11100000","00000111","00000000","00100000","00100100","00000001","10000000","00000000","00100101","00000101","11100000","10000000","00000001",
     "00100100","00100010","00100110","00100000","00101001","00101100","00101110","00000100","00000100","00000000","00000101","00000101","11110000","01010101","11010000","00011100",
     "00000101","00000101","11110000","01010101","11010000","00011100","10000100","10000100","00010100","00100000","00100100","00100100","00101001","00000101","00000001","10000000",
     "00011101","00000111","00001110","00000100","11110000","01000110","10000100","00000111","00100111","11010111","11110111","10001010","00100000","00000101","01000110","10010010",
     "10000000","01000110","10000100","00000111","00100111","11010111","11110111","10001010","00100000","00000101","01000110","10010010","00000111","00100111","11010111","11110111",
     "10001010","00000111","00100000","10000000","00000011","00000111","00001110","11111100","10000110","10010110","11010110","11110111","10000111","10010111","00100101","00101000",
     "11010111","00000110","11010111","00001000","10000101","10001000","00001111","00001110","01110111","01100110","10010111","10000111","10100111","00010111","10000111","10000110",
     "00001111","10000000","10010110","00100111","11010110","11111010","00000010","01000011","00000111","10000000","01001000","10000000","01001000","10000001","01001000","10000001",
     "10000100","01001000","10000010","01001000","10000010","01001000","10000011","10010110","01000111","10000011","10000111","10000000","11110111","10000111","10010111","11010111",
     "11010111","10001000","01110111","01111110","00010111","10000110","10000111","10010110","00001111","00100111","11010110","11111110","00000010","11110000","10010110","00100111",
     "11010110","11101010","01110100","00000110","00000101","00000101","00000000","10010110","00100111","11010110","11101000","01100000","10000000","00001000","00000110","00000101",
     "00000101","00000000","00100111","11000110","10001000","00001000","10000111","10001110","10101000","10000110","01110110","00000011","10001000","01101100","10100000","11000110",
     "10000100","10000111","10001110","10000110","00001000","00001000","00000011","01110110","10000110","11100000","01000110","10000110","10000111","10001000","10001010","00000111",
     "10000110","01110110","10011110","10100110","10000110","10101000","01000110","10000010","00000111","10000110","10000010","00001000","00001000","00000011","10000111","11110110",
     "01110111","10000110","11111010","10100110","00000111","00000111","10000110","10101010","00100000","10000101","10000000","00000110","10001010","00000110","10000110","00000110",
     "10001100","10100110","10100000","00000111","10000110","10100010","00100000","10000101","10000000","10100110","10000111","00000111","10000110","10101000","00100000","10000101",
     "10000000","10100000","11001000","10000000","10000111","10001100","10100110","10000110","11110110","00001000","00000110","01110000","00000110","10000000","10100100","00000111",
     "00100000","10000101","10000000","10100100","11000110","10001010","00000110","00000111","10010110","10000111","00000111","11110000","10100111","00000111","10101010","11000111",
     "10001010","00001000","00000111","10000110","10100110","10000111","11110111","10000110","10100110","10001010","00000111","00100000","10000101","10000000","01000111","10001000",
     "00000111","10000100","10100110","10000111","11110111","10000110","00001000","10101100","11100100","01000110","10001110","00000111","10001000","00000110","00001000","10000110",
     "11110110","01111110","10100110","10000111","00000111","10000110","10100010","11110000","01000110","10001000","10000111","10001010","10000010","00000111","11110000","11000110",
     "00000111","00000111","10000010","10000010","00000110","11110000","10100000","11000110","10001000","10000110","10000010","00000111","11110000","10100100","11000110","10001010",
     "00000111","00000110","10010010","00000111","00000111","11110000","00000111","11110000","10000111","00000111","11110000","00000111","11110000","00000111","00000111","11110000",
     "10000111","00000111","11110000","00000111","11110000","00000111","00000111","11110000","10000111","00000111","11110000","00000111","00000111","11110000","00000001","00101100",
     "00101010","00101000","00100110","00100100","00100000","00101110","00101110","00100010","10000100","11000101","00000100","00101000","00100110","10100010","10100100","10100110",
     "10101000","10101010","10101100","10101110","00101000","00101010","00101100","00101110","00100000","00100010","00100100","00100110","00001011","00001011","10001010","00001001",
     "10001001","10001110","00001010","10000101","10000101","11110000","00000111","00010101","10000101","00100111","00100111","01000111","10000111","00100000","00011010","00100110",
     "00001011","01000101","01110010","00000110","00000111","11000111","10000010","10000000","00100111","10000111","00100110","11111110","11000101","11000111","10010010","10000111",
     "00100110","11100110","01000111","00100110","00001010","10001110","10000101","10000101","11110000","00000111","00010101","10000101","00100111","00100111","01000111","10000111",
     "00100000","00011010","00100110","01110100","00000110","01000111","11000111","10001010","00000000","00100100","00000100","00100110","01100010","00000100","10001001","00100101",
     "10000101","00000100","11010000","00000101","00100101","00001001","11010000","00001001","10011110","00100000","00100100","00100100","00101001","00101001","00101010","00101010",
     "00101011","00101011","00000001","10000000","00000100","00100110","01101110","11110000","00001011","01100100","11110000","10010110","11110000","00000001","00100010","00100110",
     "11110100","00100100","00100000","00101110","00101100","00101010","00101000","00100110","00100100","00100010","00100000","01100100","00000100","00011001","00001000","10001100",
     "00011001","00000101","00001100","00001011","10011110","00000011","10001011","11011001","10000110","00001000","10011000","10000101","00000111","11010110","10000111","10000110",
     "10011111","10011000","00000100","00000110","00000110","00001000","11110000","00001111","00011010","00001010","00000101","00001110","00010011","10001000","00000110","10000111",
     "10010110","00000110","10000111","10000110","00101110","10010110","00000111","00000101","10000101","00000110","10001110","11110000","00001101","00001000","00000101","00000111",
     "00000110","00001110","00011111","00001110","00000110","00000000","00010101","10000110","01010101","00000111","10001110","10100111","00010101","01010101","10100111","00000110",
     "00000101","00000101","11011000","10010101","10000110","01010101","00000110","00000111","10010110","10000110","00001000","10000110","10001110","11110000","00000101","11010000",
     "00000101","10000011","10000101","00001000","10100000","10000111","00000110","00000110","00010111","10011000","10000111","00000110","00000111","10000110","10100000","10010010",
     "10001000","00000011","10010100","00001110","00000101","00000111","00000110","00000011","00001000","00000110","00000000","00010101","00000110","01010101","00001000","00000111",
     "01110000","00100111","00010101","01010101","10100111","10000110","00001000","00000101","11010110","10010101","00000110","01010101","00000110","00001000","00000111","01100100",
     "00000011","00001110","01101100","11010000","00000101","00001111","10001110","00001111","10000101","10001000","00000011","10100000","00001000","10000110","00000110","00000111",
     "00010111","00011110","00000111","00000110","10000111","00001000","10000110","10100000","01100000","00000011","10001000","00000101","01101110","00001111","10001110","10001111",
     "01100000","00001110","00000101","00000111","00000110","00000011","00001000","00000110","00000000","00010101","00000110","01010101","00001000","00000111","01110000","00100111",
     "00010101","01010101","10100111","10000110","00001000","00000101","11010110","10010101","00000110","01010101","00000110","00001000","00000111","01100100","00000011","00001110",
     "01101100","11010000","00000101","00000110","10001110","00001110","00000101","00100000","10000011","10001000","00001000","00000110","00010111","10010111","10000110","10001000",
     "10000111","00000011","11010111","11010111","01110111","11110111","00000111","00001000","00100000","11100110","00000101","00001110","10001110","01100100","00000110","10001100",
     "00001100","01100110","00000101","00000111","00000110","00000011","10001000","00000110","00000000","00010101","00000110","01010101","00001000","00000111","01110000","00100111",
     "00010101","01010101","10100111","10000110","00001000","00000101","11010110","10010101","00000110","01010101","00000110","00001000","00000111","01100100","00000011","10001010",
     "01101100","11010000","00000110","00000111","00000110","11010111","10000111","10000110","00000111","10011111","11100110","00000110","00001011","01101100","00100000","00100100",
     "00010101","00100100","00101001","00101001","00101010","00101010","00101011","00101011","00101100","00101100","00101101","01010101","00000001","10000000","00000101","11010000",
     "00000101","00000101","11010000","00000101","00000101","11010000","00000101","00000101","11010000","11110000","00000001","00100100","00100110","00000100","10000111","00100110",
     "00100101","00100110","00100101","11110000","00000101","00100100","00100000","00000001","11010000","00000001","00100110","00100100","00100010","00001000","00010100","00000110",
     "10000011","11110011","10000100","00000101","00010110","00000000","00000101","00000111","00000111","10010111","11101000","00000010","00001001","10010010","10000011","00000010",
     "00001110","00010100","10001111","00001111","00001000","10001110","00001110","10000101","00001000","00000110","00010111","11010111","10000011","10000101","10001000","00001000",
     "01010111","01010111","00000110","01110110","00000110","10000111","00010111","01010111","00000111","10011111","11110111","00010000","11101010","00001111","10001111","01100000",
     "10000111","10000111","00100100","11110111","10000111","10100010","10100000","10100100","10100110","00100100","00101001","00000001","10000000","10000011","00001001","00000101",
     "00000010","11110000","00001111","00001000","00001110","00011000","10001000","10011111","00000011","00000101","00000111","00000101","10011110","10001110","00000111","00000000",
     "00010101","10000111","01010101","10000111","10001110","10100110","00010101","01010101","00100111","10000101","00001000","00000101","01011000","00010101","10000111","01010101",
     "00000101","10000111","10010110","00000011","00001000","00010000","10000000","00000101","10000000","00001010","00001110","00011000","00011110","00011111","00001000","00001000",
     "00011110","00000011","10000110","00000111","10010111","00000110","10000111","00000111","00101110","00010110","10001000","10000101","00001000","00011000","10000000","00000110",
     "00001000","00010110","00010110","10000110","10010011","01010110","00000101","10011000","00001000","00000111","11010111","10000111","00000111","10011111","10011000","10000101",
     "00000110","00011110","10000000","00001000","00011110","00010101","10001110","10000011","10100000","10000111","00001000","00000101","00010111","10011000","10000111","00001000",
     "00000111","00000101","10100000","00010010","10000101","00000110","10010100","10000000","00000110","00010011","00000001","00100110","00001111","00001110","00010100","10000010",
     "10001111","00000011","10001110","10001000","10100000","10000101","00000111","00000110","10010111","10011000","10000111","10000101","00000111","00000110","10100000","00010010",
     "10001110","10001000","10010100","10000011","00001111","00001110","10000010","00010110","00100100","00000001","10000000","10000000","00000000","00010011","00000001","00100110",
     "00001111","00001110","00010100","10000010","10001111","00000011","10001110","10001000","10100000","10001000","00000110","00000101","00010111","00010111","00000110","00001000",
     "10000111","11010111","11010111","01110111","11110111","00000111","10000101","10100000","00011000","10001110","10001000","10011010","10000011","00001111","00001110","10000010",
     "00011100","00100100","00000001","10000000","10000000","00000011","00000111","01111110","01110111","10010000","10010010","01110110","01110110","10000110","00100000","00100010",
     "00100100","00100110","00000111","01100110","00010100","10000000","00000110","10010110","00000010","10000110","10000000","00000111","00000110","00000110","00000101","00000101",
     "00000100","00000100","00000011","00000011","00000010","00000010","00000001","00000001","00000000","00000000","10000000","11110101","10010110","11100101","10010110","11100101",
     "11110000","10010110","00000010","10000110","10000010","10000000","10000000","10000111","00000111","00000110","01111000","11110000","00000001","00010111","00100110","00100100",
     "00100010","00100000","00101110","00101100","00101010","00101000","00100110","00100100","00100010","00100000","00101110","11110111","00000001","00000111","10000111","00000111",
     "10000110","00100110","00000101","00000101","11100000","00000101","11000000","00011110","00000101","11000000","00011111","00000101","11000000","00010000","00000101","11000000",
     "00101100","00000101","11000000","00000010","00101110","00010111","00000111","11110111","00000111","00000111","00100010","10100111","10001110","00000111","10010100","00100111",
     "10010111","10011110","00100111","00110111","10000111","00100110","00000111","00011000","00100111","00011000","00001000","00001000","11110101","00000101","11110111","00001000",
     "11110110","00110110","00100010","10101010","00011110","11110101","10000101","10001000","00000101","00010101","01010101","00000110","01010101","11111000","00000110","00101010",
     "10011110","00011100","10011110","10011110","00010110","11110111","10000110","00010111","00000111","11110111","00000111","00000111","00100110","10010101","00100101","00100010",
     "11100000","00100111","10011010","00000111","00101100","00010111","11110100","10000111","10000100","10000111","10000100","00100111","00000100","00010111","10000111","10010111",
     "00101100","11100000","00101001","00101010","00101100","00000000","00000101","10000101","11010000","01010101","11000000","00011010","00000101","10000101","11010000","01010101",
     "11000000","00011010","00000000","00000100","00010100","11100000","11100000","11100000","00000110","00000111","11010111","00100111","10000111","10000111","00101100","00100101",
     "00000101","11000000","11100000","00010100","11110100","10000111","10000111","00000101","10000101","11100000","11100000","11100000","10000111","10000111","10000111","00001011",
     "10010101","10001011","00000101","00100010","11000000","00100111","00000101","10010101","11000000","00100111","00000101","10010101","11000000","00000101","00010101","11000000",
     "10000111","10000111","00001001","00000110","11111000","10011001","00000111","00000100","11110111","10000111","00010010","00100101","00101010","00000101","10001100","11101010",
     "11000000","00001001","00100100","00001010","00101100","10100110","00001010","00001101","10001110","00010111","10000111","11110110","10000111","10000111","00100010","00011101",
     "00000000","00100111","00000110","10010110","10000110","00000110","11010110","10001000","10000111","10010100","10100110","01010100","10011101","00011010","11011101","11011010",
     "11111100","10010100","00100111","00000100","10010100","10000100","00000100","10100110","10010110","11110110","10000110","11010110","00000010","00100111","00000110","10000101",
     "10000101","11000000","11010110","10000110","10010110","00100111","00000100","10010100","10000100","00000100","10100110","11110110","00001000","11010110","00000100","00100110",
     "00100111","10000101","10000101","11000000","11010110","10100110","00000110","10010110","11110110","10000000","00100111","00000100","00010100","10000100","00000100","01010110",
     "00010000","01010110","11110000","00100111","10010111","10010110","00100111","00000111","00011000","11110000","00010111","00000111","00000111","11110111","00000111","10010110",
     "10100101","00100010","11100000","00100111","00100000","11110111","00001110","00010111","00000111","00000111","11110111","00000111","00100010","00100111","10010111","00100101",
     "00010110","00100101","10010111","11100110","00000110","11110000","00100111","11110000","00100111","10000111","00000100","01011010","10000111","00011100","00100101","00000101",
     "10001100","11101001","01111010","11000000","00001001","00100100","00001010","11110000","00100111","00000110","10000101","10000101","11000000","01010110","10000110","10010110",
     "11010110","00010110","11110000","00000100","00000100","00101100","11000000","00100101","00000100","00100101","00000101","11000000","00100101","00000101","00000101","11000000",
     "10000101","00000101","11100000","00000101","00100101","00000101","11000000","00010100","00000101","10000101","01010100","11100000","00011000","00000101","10000101","11100000",
     "00000111","11110100","10100111","00100101","00100101","00000101","10000101","00010100","11010100","11000000","00100101","00100101","10000101","00000101","11000000","00100101",
     "00100101","10000101","00000101","11000000","00100101","00100101","10000101","00000101","11000000","00100101","10000101","00000101","11000000","00100111","11110110","10001000",
     "10100110","10000100","00010111","00000111","11110111","00000111","00000111","00000100","00101001","00100010","00011001","00010111","00100111","10000111","10010111","00000111",
     "00000111","11010110","00000101","10000101","11000000","00000100","10100111","00010100","01010100","01100100","00100111","11110110","10001000","10100110","10001010","00010111",
     "00000111","11110111","00000111","00000111","00000100","00101001","00100010","00011001","00010111","00100111","10000111","10010111","00000111","00000111","11010110","00000101",
     "10000101","11000000","00000100","10100111","00010100","01010100","01100100","00100111","11110111","10000110","10100111","10000010","00010111","00000111","11110111","00000111",
     "00000111","00000100","00101001","00100010","00011001","00010111","00100111","10000111","10010111","00000111","00000111","11010110","00000101","10000101","11000000","00000100",
     "10100111","00010100","01010100","01100100","00010111","10100111","00000111","11111001","00000111","00000100","00101010","00001001","00011001","10001110","00010111","10000111",
     "10010111","00000111","10000111","11010110","00000101","00000101","11000000","00000100","10100111","00010100","01010100","01100110","10000110","01010010","00100101","00000101",
     "11000000","00000101","11100000","00000001","00100000","00000101","00100100","00100100","00101001","00101001","00101010","00101010","00101011","00101011","00101100","00101100",
     "00101101","00101101","00000001","10000000","00000111","00101110","11110000","00010110","00000110","00000110","00000110","00001000","00100010","00101100","00000110","00000110",
     "00000000","00000110","00000101","10000110","00101000","10001110","11110000","00001000","00000011","11111000","00000110","00010110","01010110","00001000","00010011","00000011",
     "00000011","00001000","00100010","10101110","10001110","11110000","00100101","00000101","11000000","11110000","00011011","00000111","00000010","00000100","11110000","00100101",
     "00000101","11000000","11110000","00100101","00000101","11000000","00000100","11110000","10100111","00100100","10000101","00000101","10000100","11100000","11010101","00100101",
     "00000101","11000000","11110000","11110111","10000000","11110000","00100101","00011010","00000101","10001100","01001001","00111010","11000000","00001001","00100100","00001010",
     "11110000","00100101","11001010","00000101","10001100","01101001","11011010","11000000","00001001","00100100","00001010","11110000","00100101","00000101","11000000","10011001",
     "00000111","11101010","00001001","00100100","00001100","00001010","11110000","00000100","11110000","10000111","00001000","00000011","10001000","10010110","11111100","00000111",
     "01100100","00000111","01101010","01010110","00000111","11000111","00000111","00000111","01000111","00000111","00000111","00000111","00001100","10011000","01010111","00011000",
     "11101000","00010011","11010110","01010101","10010110","11010110","01010111","01110111","10000101","00010111","01101000","01111100","00001000","00000111","01100100","01101000",
     "10000101","00001000","01010111","00010011","01010011","01111000","10000110","00011000","01101000","01111110","10001000","00000111","01100110","00000111","01100100","10000111",
     "00010101","01100101","00000101","10000000","00010110","00000111","01011000","00000111","11101000","00000111","11100000","11010110","00000111","10110111","00000111","00000111",
     "01000110","10000110","00000111","10000111","10011000","10011110","10000111","11011111","11011110","00000101","01010111","01010101","01110111","00000110","00010111","01100111",
     "11111100","10000111","00000111","11100100","11100100","00000101","10000111","11010111","00010011","01010011","11110111","00001110","10010111","11100111","11111110","10000111",
     "00000110","11100110","00000111","11100100","10000111","00010101","01100101","10000000","11101000","00000111","11101010","00000111","11100000","11010111","00001000","10110111",
     "10000111","10000111","11000111","00001110","00000111","00001110","00010110","11101100","00110101","01000101","00000101","10000000","00000101","00000101","10000000","00000111",
     "11110000","11010111","00001000","11110000","00000111","10000110","01111110","11010110","00000111","11110000","00000111","00000110","01110010","01010110","00000111","11110000",
     "10011000","11010110","11011111","01011110","10010111","01010110","11100111","10011110","11011110","00010011","01010101","01110110","10000111","10010110","11100110","11111110",
     "10000110","00000110","11101110","11111100","00001110","10000110","10000110","11010110","00010111","11010111","11110110","10000101","10010111","01100111","01111110","00000111",
     "00000111","01101000","01110110","00000110","00000111","00010101","00000111","11100101","11110000","01010111","10010110","11100110","11010011","11011111","01010111","10011110",
     "11011110","10011000","01010111","01101000","01011000","00010110","01110011","10000101","00010011","01101000","11111110","10001000","10000111","11100100","11110010","10000111",
     "10001000","10001000","11010111","00011000","01011000","11111000","10000011","10011000","11100101","11111110","10000101","00001000","11101110","11111100","00000111","10000101",
     "10010111","00001111","11100111","00000111","11110110","11011000","01110111","01010110","10001110","10000101","10000110","11011000","10000111","10000110","00000110","10000110",
     "11110100","00000110","11011000","10000110","11101010","10001000","10000101","00000101","10000000","00000111","00000111","11110110","10010110","11111110","00010101","10000110",
     "01111100","10000101","00000101","10000000","11010111","00001000","11110000","01010110","00000111","11110000","11010110","00000111","11110000","00000101","00000101","10000000",
     "10000111","00001000","11110000","00000111","11110000","10000110","11110000","00000111","11110000","00001110","11110000","00000101","00001000","11110000","00000101","10000111",
     "11110000","11000111","11110111","00001000","10010010","00000111","11111110","01110111","00000111","10011000","11110110","00000111","01101100","01111100","10000110","00000111",
     "10101000","10000111","10000110","10101110","11101000","00000111","10000111","11110111","10000111","00000111","10000101","01101000","10000000","00000111","01111100","11000111",
     "00000111","10000101","00001111","01101000","10000000","11000110","00000111","01110111","00001111","10000101","10000000","11000110","00000111","01110111","00001111","10000101",
     "10011010","11110000","10100110","10100010","10101111","10101111","10101110","10101110","10100011","10101000","10000101","00100000","10100110","00100010","00100100","00100110",
     "00101000","00101010","00101100","00101110","00000111","00101110","01101000","11110000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
  signal ram_symbol2 : ram_type := (
     "00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","00010001","01010001","01100001","01110001","10100001","10110001","11000001","11010001",
     "11100001","11110001","00000001","00010001","11000001","11010001","11100001","11110001","00000001","01010000","11000001","10000001","01000001","00000001","11000001","10000001",
     "01000001","00000001","11000001","10000001","01000001","00000001","11000001","10000001","01000001","00000001","00000001","00100000","00000000","10000001","00000000","10000001",
     "00000000","00000101","00000001","10110101","00000101","01000101","01011111","00000000","01000101","11000001","00000000","10000101","10110101","00000101","01000101","10100001",
     "00000110","00000001","00011111","01000001","00000000","00000101","01000101","00000000","10000101","00000101","10010000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00110010","00110110","01100001","01100101","01101001","01101101","01110001","01110101","01111001",
     "00000000","00110010","00110110","01000001","01000101","01001001","01001101","01010001","01010101","01011001","00000000","01010101","00000000","01111000","01100011","01010000",
     "01100101","01110010","01101110","01100111","00100000","01001000","00000000","01111000","01100011","01000101","01110101","01100111","01110010","01110010","00100101","01110100",
     "01110100","01110011","01010100","00100000","00100000","01100101","01101101","01101001","00101110","00000000","01000101","00110011","01000001","01110010","01110010","00100000",
     "01100010","00100000","01111001","01101111","01101000","01101110","01100101","01100001","00001010","00000000","01100001","01010100","00100000","00000000","00100000","01100110",
     "01100001","00100000","00100000","01100001","01100101","01100110","01100011","01101101","00101110","00000000","00100000","01101001","01101001","01110010","01110000","01101101",
     "01110010","01101111","01101111","01100001","00001010","01101111","01100101","01101110","01110100","00100000","00100000","01100001","01100101","01100110","01100011","01101101",
     "00101110","00000000","00100000","01100110","01100001","00100000","00100000","01100001","01100101","01100110","01100011","01101101","00101110","00000000","00100000","01101001",
     "01101001","01110010","01110000","01101101","01110010","01101111","01101111","01100001","00001010","01110101","01010010","00100000","01110100","01100011","00100101","00100000",
     "01101000","01100100","00100000","00110000","00000000","01110101","01010010","00100000","01110010","01100011","00110000","00110100","00100000","01110101","01100010","01111000",
     "01111000","00000000","01110101","01010010","00100000","01110100","01110010","01111000","01111000","01110011","01101100","01100101","00100101","00001010","01110010","01110010",
     "01101001","00100000","00100000","00001010","01110100","01110100","01110011","00100000","00100000","00001010","01110100","01110100","00100000","01100011","00100000","00000000",
     "01100101","01101001","00101111","00100000","00100000","00000000","01010010","00100000","01110100","01100101","01100101","01110010","00100000","01110011","00110000","01100011",
     "01101111","00100000","01101001","01100101","01110100","00000000","01100101","01101001","00100000","00100000","00100000","00001010","01000011","00101110","00000000","01101101",
     "01100101","01100101","01101111","00100000","00000000","00100000","01100001","00101100","01100101","01101011","01101100","00000000","01101101","01100101","01101100","00100000",
     "00100000","00000000","01000001","00000000","01101101","00100000","01100001","01101110","00100000","00000000","01100101","01100011","00100000","00100000","00100000","00110000",
     "00000000","01100100","01100011","01110100","00100000","00111010","00100101","00001010","01100100","01100011","01110010","00100000","00111010","00100101","00001010","01100100",
     "01100011","01110100","00100000","00111010","00100101","00001010","01100100","01100011","01100001","00100000","00111010","00100101","00001010","01110010","01110100","01100101",
     "01101001","01110110","01100100","01100100","01100101","01000101","01000101","00100000","00100000","00100000","00100000","01101111","01101110","01110101","00101110","00000000",
     "01110010","00100000","01100101","01100100","00000000","01101110","00100000","01101001","01100101","01100101","01101001","01100110","01110100","01100101","01100101","01100001",
     "01110011","01101100","01100101","01101101","01100101","01110100","01100101","01110100","01101110","01101011","01101110","01100001","01110010","00000000","01100001","00000000",
     "01100001","00000000","01100001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00101110","00110001","00000000","00101110","01010100","00000000","00110011",
     "00110100","00000000","00101110","01010100","00000000","00110101","00101011","00000000","00110001","00101101","00000000","00110111","00110011","00000000","00101110","00110001",
     "00000000","00101110","00110000","00000000","00110010","00110000","00000000","00110001","00110000","00000000","00101110","00110000","00000000","00110001","00000000","00110011",
     "00000000","00110111","00000000","00110010","00000000","00000010","00000011","00000100","00000100","00000101","00000101","00000101","00000101","00000110","00000110","00000110",
     "00000110","00000110","00000110","00000110","00000110","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",
     "00000111","00000111","00000111","00000111","00000111","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","01010000","10100111","00000000","00000111","00100101","11110101","00000101","00000111","00000000","10000111","00000000","11000001","00000000","10000001",
     "00000000","00000000","11000111","00000000","01000001","00000000","00000000","00000000","10110101","00010110","00010101","00010101","00000110","11111111","00010110","11010111",
     "00000111","00000111","11100111","00010111","00100101","00010111","00000111","11111111","00010111","11100111","00000111","00000111","11010111","00010110","00110101","00010111",
     "00000110","11111111","00010110","11010111","00000111","00000111","11100111","00010111","01000101","00010111","00000111","11111111","00010111","11100111","00000111","00000111",
     "11010111","00010110","01010101","00010111","00000110","11111111","00010110","11010111","00000111","00000111","11100111","00010111","01100101","00010111","00000111","11111111",
     "00010111","11100111","00000111","00000111","11010111","00010110","01110101","00010111","00000110","11111111","00010110","11010111","00000111","00000111","00010111","00010111",
     "11100110","11111111","00010111","11110101","00000111","00000101","00000000","10100101","11110101","00010110","00010110","00010101","00000110","11111111","00010110","11000111",
     "00000111","00000111","11100111","00010111","00010111","00100110","00000110","11111111","00010110","11000111","00000111","00000111","11100111","00010111","00110110","00010111",
     "00000111","11111111","00010111","11100111","00000111","00000111","11000111","00010110","01000110","00010111","00000110","11111111","00010110","11000111","00000111","00000111",
     "11100111","00010111","01010110","00010111","00000111","11111111","00010111","11100111","00000111","00000111","11000111","00010110","01100110","00010111","00000110","11111111",
     "00010110","11000111","00000111","00000111","11100111","00010111","01110110","00010111","00000111","11111111","00010111","11100111","00000111","00000111","00010111","00010111",
     "11010111","11111111","00010111","11100111","00000111","00000111","10000101","10100111","11110101","00010110","00010111","00010111","00000110","11111111","00010111","11110101",
     "00000101","00000101","10100110","00010110","00100111","00010101","00000110","11111111","00010110","11010101","00000101","00000101","11110101","00010111","00110111","00010101",
     "00000111","11111111","00010111","11110101","00000101","00000101","11010101","00010110","01000111","00010101","00000110","11111111","00010110","11010101","00000101","00000101",
     "11110101","00010111","01010111","00010101","00000111","11111111","00010111","11110101","00000101","00000101","11010101","00010110","01100111","00010101","00000110","11111111",
     "00010110","11010101","00000101","00000101","11110101","00010111","01110111","00010101","00000111","11111111","00010111","11110101","00000101","00000101","00010101","00010101",
     "11100111","11111111","00010111","11110101","00000101","00000101","00000000","10100101","11110101","00000101","00011000","00000111","00010110","00010101","00001000","11111111",
     "00010101","10110111","00000111","00000111","11000111","00010110","00010111","00100110","00000101","11111111","00010101","10110111","00000111","00000111","11000111","00010110",
     "00110110","00010111","00000110","11111111","00010110","11000111","00000111","00000111","10110111","00010101","01000110","00010111","00000101","11111111","00010101","10110111",
     "00000111","00000111","11000111","00010110","01010110","00010111","00000110","11111111","00010110","11000111","00000111","00000111","10110111","00010101","01100110","00010111",
     "00000101","11111111","00010101","10110111","00000111","00000111","11000111","00010110","01110110","00010111","00000110","11111111","00010110","11000111","00000111","00000111",
     "00010111","00010111","11010110","11111111","00010110","11010111","00000111","00000111","10000111","11100111","00010110","11110111","00010111","00010111","00000110","11111111",
     "00010110","11010111","00000111","00000111","11000111","00010110","00100111","00010111","00000110","11111111","00010110","11000111","00000111","00000111","11010111","00010110",
     "00110111","00010111","00000110","11111111","00010110","11010111","00000111","00000111","11000111","00010110","01000111","00010111","00000110","11111111","00010110","11000111",
     "00000111","00000111","11010111","00010110","01010111","00010111","00000110","11111111","00010110","11010111","00000111","00000111","11000111","00010110","01100111","00010111",
     "00000110","11111111","00010110","11000111","00000111","00000111","11010111","00010110","01110111","00010111","00000110","11111111","00010110","11010111","00000111","00000111",
     "00010111","00010111","11100110","11111111","00010111","11100111","00000111","00000111","00000101","10100111","11110101","00000101","00010101","00000110","00010111","00010111",
     "00000101","11111111","00010111","11110101","00000101","00000101","11000101","00010110","00100111","00010101","00000110","11111111","00010110","11000101","00000101","00000101",
     "11110101","00010111","00110111","00010101","00000111","11111111","00010111","11110101","00000101","00000101","11000101","00010110","01000111","00010101","00000110","11111111",
     "00010110","11000101","00000101","00000101","11110101","00010111","01010111","00010101","00000111","11111111","00010111","11110101","00000101","00000101","11000101","00010110",
     "01100111","00010101","00000110","11111111","00010110","11000101","00000101","00000101","11110101","00010111","01110111","00010101","00000111","11111111","00010111","11110101",
     "00000101","00000101","00010101","00010101","11100111","11111111","00010111","11110101","00000101","00000101","10000110","11110101","00010111","11110111","00010111","00010101",
     "00000111","11111111","00010111","11100101","00000101","00000101","11010101","00010110","00100111","00010101","00000110","11111111","00010110","11010101","00000101","00000101",
     "10100111","00010111","00110111","00010101","00000111","11111111","00010111","11100101","00000101","00000101","10100110","00010110","01000111","00010101","00000110","11111111",
     "00010110","11010101","00000101","00000101","10100111","00010111","01010111","00010101","00000111","11111111","00010111","11100101","00000101","00000101","10100110","00010110",
     "01100111","00010101","00000110","11111111","00010110","11010101","00000101","00000101","10100111","00010111","01110111","00010101","00000111","11111111","00010111","11100101",
     "00000101","00000101","00010101","00010101","11110111","11111111","00010111","11110101","00000101","00000101","00000000","10100101","11110101","00000101","00010110","00000111",
     "00010111","00010101","00000110","11111111","00010101","10110101","00000101","00000101","11010101","00010110","00010101","00100111","00000110","11111111","00010101","10110101",
     "00000101","00000101","11010101","00010110","00110111","00010101","00000110","11111111","00010110","11010101","00000101","00000101","11000101","00010110","01000111","00010101",
     "00000110","11111111","00010110","11000101","00000101","00000101","11010101","00010110","01010111","00010101","00000110","11111111","00010110","11010101","00000101","00000101",
     "11000101","00010110","01100111","00010101","00000110","11111111","00010110","11000101","00000101","00000101","11010101","00010110","01110111","00010101","00000110","11111111",
     "00010110","11010101","00000101","00000101","00010101","00010101","11100110","11111111","00010111","11100101","00000101","00000101","10000111","11110101","00010111","11110111",
     "00010111","00010101","00000111","11111111","00010111","11100101","00000101","00000101","10100110","00010110","00100111","00010101","00000110","11111111","00010110","11010101",
     "00000101","00000101","11100101","00010111","00110111","00010101","00000111","11111111","00010111","11100101","00000101","00000101","11010101","00010110","01000111","00010101",
     "00000110","11111111","00010110","11010101","00000101","00000101","11100101","00010111","01010111","00010101","00000111","11111111","00010111","11100101","00000101","00000101",
     "11010101","00010110","01100111","00010101","00000110","11111111","00010110","11010101","00000101","00000101","11100101","00010111","01110111","00010101","00000111","11111111",
     "00010111","11100101","00000101","00000101","00010101","00010101","11110111","11111111","00010111","11110101","00000101","00000101","00000000","00000000","00000000","00000001",
     "10010001","01000001","00010001","10000001","00100001","00110001","01010001","01100001","01110001","10000001","10010001","10100001","10110001","00000111","00000101","00000110",
     "00001000","00000000","01001000","00000111","00001101","00010111","00010111","00000000","00000110","00100111","00000111","00000110","00000101","01000111","00000110","10000111",
     "00000000","00000111","11110110","00000000","00001101","00000000","11111010","10001010","00010111","11110110","00000101","00000000","11110001","00000000","00010000","00010000",
     "11000001","00001100","11101100","00000111","01010110","11111011","00001110","01100000","00001011","00000100","00000000","01100001","01010000","11000001","01100100","11100000",
     "11110000","00000011","01100100","00010100","00001101","10000000","11111010","00000000","11111010","00001101","01100000","11111011","11111010","01001011","00011010","11111011",
     "00000100","00001101","00001100","01001011","01010000","10100100","11111011","01011100","10011010","00000100","00001010","00000000","01010000","01010100","00100100","00000100",
     "00010000","00010111","00000110","11100101","00100111","10110111","11110100","11110110","11110000","00110100","01100000","11111011","11110111","11111011","00010100","00000100",
     "00000100","00000000","11010000","10000100","11000001","10000001","00000100","00000001","01000001","11000001","10000001","01000001","00000001","11000001","10000001","01000001",
     "00000001","11000001","00000001","00000000","11100111","00001101","00100111","00000000","00000111","00000110","10011111","00000000","11001000","10011111","00000000","01011111",
     "10110000","11110110","11010000","00001101","00000000","11000001","10000000","00001001","01000101","00011001","00110100","00000101","00001001","11111000","00000111","01000101",
     "11111000","01000101","11011111","11110110","10110000","11011111","00000000","11110100","10000000","11110100","00100100","10011111","11100110","01011111","00000000","11110100",
     "00010100","00011111","00001011","11111011","11011111","11101011","00001011","00000111","01011111","10100000","11110101","00000001","01000111","00000111","11110111","00000111",
     "10100111","00000000","00000001","01000111","00000111","11110111","00000111","11010000","11110111","10011111","00000001","10000001","00010001","10000001","10010001","00100001",
     "00110001","01000001","01010001","01100001","01110001","10010001","10100001","10110001","10110001","11000001","11010001","11100001","11110001","00000001","00010001","00000101",
     "01000001","10000001","00000111","00000001","00000000","00000000","00000000","00000101","00001001","10001011","11001010","11001001","00000000","01010000","11100111","11111011",
     "00010100","00011011","00010100","00000111","00001011","00000001","00000110","00010000","10100000","00000001","11010000","00100110","10110110","01000111","00000111","11110111",
     "00000111","11001001","11010111","00011001","00001001","00000110","11000001","10000001","01000001","00000001","11000001","10000001","01000001","00000001","11000001","10000001",
     "01000001","00000001","11000001","00000001","00000000","01000111","00000111","11110111","00000111","00000111","11011111","00010100","00000000","00000000","00000101","11110111",
     "00010100","11100110","00100111","01110111","00000111","00000111","00010111","00000100","00010100","00010100","00000101","11110111","11100110","00000101","11110111","10010000",
     "11100110","10100000","11110000","11100101","11100000","11110000","11000101","11110101","11000000","10100110","11110101","11110110","01110000","11000101","00100110","01000110",
     "00000110","00000110","00000111","00000100","00011111","01000111","00000100","01011111","00000111","00000100","10011111","10000111","00000100","11011111","00010100","01110000",
     "00010100","11111000","11110110","11000101","00000000","00100110","11000101","10100110","00000110","00000110","00010100","10010000","00010100","00000101","11110111","11100110",
     "10100000","11100101","00000101","00000000","11011111","00000000","10010000","00100110","11010111","00010100","00010110","10110110","00000100","00000110","00000101","11110111",
     "11100110","11011111","00001100","00100100","00100100","01001100","00000110","11010000","00000111","11011111","00000100","00000111","00000000","01001100","00001100","00000101",
     "00001011","10011111","00011100","00000101","00011100","00000111","10011111","00000100","10100000","00011111","00000100","00001100","01001100","00000100","00000100","00000110",
     "00000111","00000100","11000000","11100110","10000101","00010110","00000110","00000101","00000111","10000110","00000111","10010000","01000100","01001011","11101011","11000100",
     "11110100","00010111","00010110","10010111","11000111","00010111","11100111","00000111","10001011","00110111","00000111","11000100","00000100","00001011","10000101","00000111",
     "01000111","01000111","11000111","11110101","11000100","11110100","11111011","10011011","10010111","00000100","00010111","10100110","10010101","00010100","00100111","10110110",
     "10010111","00100100","11110110","00000111","00011100","11010100","10010110","00001011","00000100","00000000","11010000","10011011","00011100","00000111","10011111","00000100",
     "11110000","11000110","00001100","00000000","01001100","11011111","00000100","10000000","01011111","00000100","00000111","11110110","00000111","00001100","00011011","01001100",
     "11111011","00011100","10010000","00000100","00000000","00000111","11010000","00011100","10010101","00000111","10011111","00000101","00000100","01010000","00011011","11111000",
     "11111011","00001100","00001000","00000111","00001011","00000001","00000110","00000000","10011111","00000000","10010000","00100111","11100110","00010101","00010111","10110111",
     "00000101","00000111","00000101","11110110","11001000","00000101","01011111","00001100","00100100","01001100","11110111","11110110","11000111","00100100","01011111","11000000",
     "00100111","01001100","10100000","00000101","01000000","11000000","00001100","00000111","01001100","11000101","00000000","01000110","00000111","00010111","00100111","00110111",
     "01000111","01010111","01001000","01000101","01001110","01000011","01001000","11111000","11110101","11111110","11110011","11111000","01000101","00000110","10100110","01110110",
     "01010110","11110110","11000110","11100110","01100110","11010110","00010110","00001000","00000101","00000011","00000010","00001111","00001110","00001111","00000011","00001110",
     "00001000","11100110","00000101","10100000","11110101","10000001","11100001","11100001","11100001","11100001","11100001","01110001","01010001","10010001","11110001","11000001",
     "11100001","01100001","11010001","00000001","10110110","10100001","00000111","00000111","11110110","11100001","00000111","00010000","11010111","11110110","00000100","00000000",
     "00001011","11010001","11000000","00010000","10000001","10001011","11000000","11000001","11011011","00100100","00100100","00000111","00000111","11011111","11000000","00001100",
     "01001100","11000101","00001001","01011111","00000100","00000000","11011111","00001100","01001100","00000111","00000110","00110000","11000101","01000000","10100110","10100000",
     "01000000","00110000","00100000","10100110","00001000","11001001","00000110","11000001","10101001","00000110","00001000","10100001","11001001","00000110","00000001","01100101",
     "11000011","00000001","00010111","10000101","11100000","00000101","00000110","00110000","11001000","01000000","10100000","00000001","10111110","00110100","00000110","00000110",
     "00010011","11001001","00000110","11001110","00001001","00000110","00010011","00000101","11001001","00000110","00000001","10110110","00010101","10100110","00000001","00100111",
     "10000101","11100000","10110101","00010100","00000110","00110000","11001000","01000000","10100000","00000001","10111110","00110100","00000110","00000110","00010011","11001001",
     "00000110","11001110","00001001","00000110","00010011","00000101","11001001","00000110","00000001","10110110","00010101","10100110","00110111","00000001","10000110","11100000",
     "11000101","00010100","00000111","00110000","11100101","01000000","10100000","00000001","11000011","00110100","10100111","10100111","00001000","11101001","00000111","11100011",
     "10101001","00000111","00001000","10100101","11101001","00000111","00000001","11000111","00010110","10110111","00000111","11110110","00000111","11010100","10000110","00001011",
     "00001101","00000000","11010001","10000000","11000001","10101011","11010100","10010110","11110110","00001011","00000100","10000001","11010001","00000000","11000001","10001011",
     "00000111","11010100","00000000","00010000","00011011","01100110","10010111","11001011","11110111","11110100","00010100","00010100","00000111","11001111","00100111","01001100",
     "00000100","00001100","10100000","00000101","00011111","00001100","00000111","01001100","01011111","00101011","00000111","00000111","00001011","00011100","00011100","00000111",
     "00000111","11001111","00010111","10000000","10011111","10010000","00000100","00001011","00000000","10011011","11000000","11110000","01011111","11001010","10011111","11110110",
     "11010100","10010110","00001011","00001101","00000000","11010001","11000000","11000001","10111011","11010100","10100110","00011111","00000000","11000001","00010000","00000001",
     "00010111","10000101","11100000","00000101","00100000","00000110","00000001","10110110","00000000","10110110","00100100","00000001","00100111","10000101","11100000","10110101",
     "00010100","00000110","00000001","10110110","00000000","10110110","00100100","00000001","00110111","10000110","11100000","11000101","00010100","00000111","00000001","11000111",
     "00000000","00100100","11000111","11011111","11100110","00000100","00000111","00010000","10000001","00001011","11010001","10000000","11000001","00010000","00011011","11011100",
     "00000000","00100000","00010000","00010111","11100110","11111011","10110111","10000111","11110110","00011111","00000001","00001001","00001111","00001100","11011111","10010000",
     "11000101","10100000","00000110","00000001","10111000","00100100","10101001","00000101","00000110","10101000","00011111","10010000","11000101","10100000","00000110","00000001",
     "10111000","00100100","10101001","00000101","00000110","10101000","10011111","10010000","11100101","10100000","10100111","00000001","11001000","00100100","10111001","00000101",
     "10100111","10111000","10011111","10010000","11000101","10100000","00000110","00110000","00100000","00010000","10101001","00000101","00000110","10100001","10011111","00100000",
     "00010000","00000000","10011111","00000111","00000100","00000000","10011111","00001100","00011011","01001100","11111011","00011100","00011100","00000111","00000111","01001111",
     "00001101","10001111","10011011","00010100","11110100","00011011","11111011","11101011","11001111","11100110","00001100","00000111","01011111","00000001","00100001","00010001",
     "10000001","10010001","00110001","00000101","01110100","00010111","11110100","00000111","00000101","00110100","11110101","01000101","01110100","10110111","00000101","10000100",
     "00000111","00010000","11010111","00000100","00000101","00000100","00000111","11111001","00000100","10001111","10001001","10100100","00000100","10001001","11000001","10000001",
     "00001001","01000001","00000001","11000001","00000001","00000000","00100000","00000101","11010101","00100000","00100100","00000100","01000100","10000100","11110111","11000000",
     "11100100","00000101","00001001","00000111","10100100","10000100","00011111","00000111","10000100","01010000","11000100","00000101","00001001","00000111","10000100","10100100",
     "10011111","00000001","10010001","00100001","01000001","00010001","10000001","00110001","00000101","00000101","00000110","01110100","00010111","11110100","00000111","00110100",
     "11110101","01000101","01110100","11110101","00000101","10000110","00000111","00010000","11010111","00000100","00000101","00000100","00000111","11111010","00000100","00001111",
     "10001010","10100100","00000100","10001001","00001001","01110100","00010111","11110100","00000111","00110100","11110101","01000101","01110100","11110101","10000100","00000111",
     "00010000","11010111","00000100","00000101","00000100","00000111","11111001","00000100","11001111","10001001","10100100","00000100","10001001","11000001","10000001","00111010",
     "01000001","00000001","11000001","10000001","00000001","00000000","00100000","00000101","11010101","00100000","00100100","00000100","01000100","10000100","11110111","11000000",
     "11100100","00000101","00001010","00000111","10100100","10000100","10011111","00100000","00000101","11010101","00100000","00100100","00000100","01000100","10000100","11110111",
     "10000000","11100100","00000101","00001001","00000111","10100100","10000100","10011111","00000111","10000100","00010000","11000100","00000101","00001010","00000111","10000100",
     "10100100","11011111","00000111","10000100","10010000","11000100","00000101","00001001","00000111","10000100","10100100","10011111","00000110","00100101","00100101","11110101",
     "00000000","00000101","00000111","00000111","10000111","00000111","11100111","11110101","00000101","00000111","00000111","10000111","00000111","11100111","11110101","00100101",
     "00100101","11110101","00000000","00000101","11110101","00100101","11110101","00000000","00000001","10000001","00010001","10000001","10010001","00100001","00110001","01000001",
     "01010001","01100001","01110001","10010001","10100001","10110001","01000101","00000001","00000101","01000101","00010000","10110001","00000000","00000000","00000000","00000000",
     "11000001","11110110","11010001","00000111","00000100","01000100","00000111","00000100","00100111","11010111","11000000","01000111","11000001","00100111","11010111","00000111",
     "00000111","00000000","11000000","00000100","00000111","00000100","11010100","00000111","00000111","01000111","00010101","00000101","00000111","00000101","00010111","00000110",
     "10010111","00010111","11101000","00000111","00001000","00000111","00000110","00000110","11100111","00000100","11110110","11010100","11000001","00000111","00010111","00001011",
     "00000111","11110001","00010110","00000110","00000110","11001000","00100101","11000111","11111000","00000111","00000111","11110001","10110000","00000100","00000100","00000111",
     "01000111","01001001","11010111","11101001","00000111","00000111","11100111","11000001","00001001","00000111","01000100","11000001","00100111","11100111","00000100","00000100",
     "00000100","00000100","01000100","11000001","00000111","10011111","00000100","10100001","00000100","00000100","01000100","01001001","00010000","11111001","00000100","11100100",
     "00000000","11111001","00100100","00000000","00000000","00010000","00011110","00000100","00000000","00000110","00010111","00000110","11110011","00000011","00000100","00000011",
     "00000110","00000111","00000110","00000100","01000111","01000100","00000101","00000110","00001000","10001000","00000110","00000110","11010101","00000101","00100101","00000110",
     "00001000","00000110","10001000","00000110","11010101","00100101","11010110","11010000","00000100","00000100","11110110","00001000","11011000","00000110","00000111","00000110",
     "00000100","00000100","11110110","00000100","00001000","00000110","00000110","11011111","01000100","01000001","00000111","11100111","00000100","00000100","00000100","00000100",
     "10011111","00000111","11110111","00000111","11011111","00000100","00001000","11101110","00010011","00000100","00000100","00000000","00000000","00000000","00011111","00000100",
     "01000100","00000100","00000111","11100110","01011111","01000111","01000001","00000111","11010111","00000111","00000111","10011111","01000110","00011110","00000111","00010111",
     "00001110","00010111","11101000","00000111","00001000","11011111","00000100","00000100","01000100","11000001","00000111","00001111","00000100","10100001","00000100","11000001",
     "10000001","01000001","00000001","11000001","10000001","01000001","00000001","11000001","10000001","01000001","00000001","11000001","00000001","00000000","10110001","00000001",
     "10110000","00000100","00010000","11110001","10001100","11110001","00000100","00000000","00000000","00000001","00010000","00000001","00001101","00000000","00010111","11110001",
     "00001101","00011011","00001101","10000001","11111011","10000001","00001011","00001100","00001101","01001101","01001101","00001010","00000100","11110100","00000111","00110100",
     "11110101","01000101","01110100","11110101","10001100","00000111","01000111","00000100","00000101","00000100","00000111","00011111","11111011","00000100","00011011","10101100",
     "00001000","00011010","00001001","00001010","11111010","00000111","00111010","11110101","01000101","01111010","11110101","10001100","00000111","01000111","00001010","00000101",
     "00001010","00000111","01011111","11110100","00001010","00010100","10101100","00001000","00011001","10011011","10010000","00001101","00001101","11111100","00001001","11111001",
     "00000111","00001011","00001100","00001101","00001101","11111100","00001101","00001001","00000111","00000111","11011111","00001101","11111011","00001101","00011111","00001101",
     "00001101","00000001","00001001","00010000","11110111","10000001","00010111","11110001","00000100","00000000","00010000","10000001","00000111","01000000","11001100","00000101",
     "00000100","00000111","10001100","10101100","01011111","00100000","00000101","11010101","00100000","00101100","00001100","01001100","10001100","11110111","00010000","11101100",
     "00000101","00000100","00000111","10101100","10001100","00011111","10000001","00000111","10000000","11001100","00000101","00001011","00000111","10001100","10101100","11011111",
     "00100000","00000101","11010101","00100000","00101100","00001100","01001100","10001100","11110111","01010000","11101100","00000101","00001011","00000111","10101100","10001100",
     "10011111","11000001","01011111","00000000","00010000","01000000","11110101","00000101","11111111","00000111","00000101","10000101","11100101","00110101","11100101","11100101",
     "00001111","01000101","00100101","11111111","00000111","01001111","11100110","10001111","00000101","11111000","11100101","00010101","01100101","11110000","11110111","11101111",
     "11111111","00000101","00000101","00000110","11111111","00000011","00000000","11110010","10000110","11101110","01001000","11111110","00001000","00000011","01110011","00110111",
     "10000111","01110011","11100110","01100111","11010101","10000111","00000110","11110111","11111000","01011000","00000101","00001110","00001110","00011000","00010101","00000111",
     "00000111","01010000","11110101","00000000","00010000","11110011","01000111","10100110","11011000","00000111","00010110","00000111","00000111","00010000","00010000","00000101",
     "00000000","00000000","00000000","00011111","00000111","00000000","00000101","00010111","00000101","11110111","00000111","00001111","00000101","00000111","00000110","00000111",
     "01000110","01000111","00000011","00001000","00000101","10000101","00001000","10101000","00000011","00001110","00101110","00001000","00001110","00001000","10001110","11011000",
     "00001110","00100011","01010101","10100000","00000111","00000111","11110110","00001000","00001000","00001000","00000111","00000110","00000111","00000111","11110110","00000111",
     "00001000","00001000","00001000","11011111","00000110","11110111","00000110","00011111","00000111","00001000","01111111","00011111","00000101","00000000","00010000","00000110",
     "00001000","00011000","10000111","00000111","11001000","00000111","01100111","11111000","00000111","00010110","00000111","00000111","01011111","00000101","00000000","00000101",
     "00000011","00001000","00011111","00000011","00001000","01011111","00000110","10001000","11101000","00000110","01000111","11110111","00010110","00000101","11111000","00000101",
     "00000110","00001000","11111000","01000111","11110110","00000101","01001000","11100111","00100101","11100111","00000000","00000000","00001000","00000000","00000101","01000101",
     "00000101","01000111","00000111","11000111","11010111","00000111","00000110","11010111","00000111","00000000","01000101","01000101","11100101","00000101","11010101","11100101",
     "10100101","00000000","00100101","00000111","00000101","01000101","00100111","11100111","00000000","01000101","00100111","11100111","00000101","00000101","00000000","00000101",
     "01000101","00000101","00000111","11100111","01000000","01000101","00000111","11100111","00000101","00000101","00011111","00000000","00000000","00000000","00000101","00000000",
     "10000000","00000111","00000101","11100101","00000101","00000111","00000000","00000101","00000001","01010001","01100001","01110001","10000001","10100001","00010001","10000001",
     "10010001","00100001","00110001","01000001","10010001","00000101","00000101","00000110","00010000","00010000","00001011","00000000","00000000","00000000","00011100","00001010",
     "00000000","00000100","00010100","00000100","01010100","00001010","00000100","00001001","00000100","01000100","01001010","00001100","00001011","10100000","00000100","00000100",
     "11111001","00001001","11111001","00000111","00000100","00001001","00000100","00000100","11111001","00000100","00001001","00000111","00000111","11011111","00001010","11110100",
     "00001010","00011111","00000100","00000100","00001001","10101100","00011010","00001011","00000000","00010000","11000001","10000001","00001011","01000001","00000001","11000001",
     "10000001","01000001","00000001","11000001","10000001","01000001","00000001","00000001","00000000","00000000","00010000","00000000","00000000","00000000","00000000","00000000",
     "00000000","11010111","11000111","00000010","00000111","00001111","00000111","00000001","00000110","11010111","11110111","11010111","00100111","11100111","00000000","00000010",
     "10000111","00000000","00000111","11100111","00000000","00000000","00000000","10000111","00000111","11000111","01000111","10100101","10100101","11100111","10110111","00000000",
     "00000001","01000000","00000000","00010001","01010000","11000001","00000001","00000000","00000001","10000001","00000101","00000000","01000000","01000101","00010001","11001111",
     "00000000","00000000","11000101","11001111","00010000","11110100","11000001","10000001","00000001","00000000","00000101","00000000","10000101","01001111","00000000","00000001",
     "10000001","10010001","00010001","00100001","11000101","00000101","00000101","00000101","00000000","00001001","00010000","00000100","00001111","10000100","01001111","10100100",
     "11110000","00000100","10001111","10000100","11001111","10100100","00000100","00010100","10011001","11000001","10000001","01000001","00000001","00000000","00000001","00000000",
     "10100100","00010000","11111001","00010000","10011111","00000101","00000110","00000001","01000111","00000111","11110111","00000111","11010111","00010101","00000101","00000110",
     "00000000","00000101","00000110","00000001","01000111","00000111","11110111","00000111","11010111","00010101","00000101","00000110","00000001","01000111","00000111","11110111",
     "00000111","10100000","11110111","00000000","11110101","00010000","00000110","01100111","00010101","00000110","00000110","01110110","11010111","00000111","00000000","00000000",
     "00110110","01000000","00000111","00000000","01000101","00001000","10000000","11000000","00110111","11110110","00100111","00010111","00000111","00100111","11100101","00010110",
     "10011000","00000111","00000110","00000111","00000110","01101111","10000000","00000111","00001110","01110111","00010111","00000111","00100111","00000111","00110111","00000111",
     "11000010","01000111","00000111","01010111","00000111","01100111","00000111","11100010","01110111","11100111","01010111","11010111","01110110","11010111","00000111","00110110",
     "00000111","00001111","00110111","11110110","00100111","00010110","11100101","00000110","01011000","00000111","00000110","01101111","01000000","10011111","00000110","00000111",
     "00000110","01101111","10101000","00000101","00000000","00001110","11010000","00000110","00000111","00000110","01101111","10101000","00000000","00000000","00000101","00000000",
     "00001110","00010000","00000101","00000111","00000110","11000000","00010111","00000110","00000101","00000110","11110110","10010000","00011000","11000011","00010101","00010111",
     "00000110","00100111","00000110","00000110","11100000","10010000","11000000","11110110","00000110","11001000","00010111","00010111","00000111","00000110","01100110","00000110",
     "00000110","11110110","00000110","00000101","00010110","11010101","00010111","00000110","11000000","00010111","11100110","01010000","10010000","11000000","00000110","11110110",
     "11110111","00000110","11101000","01000101","00000110","00010000","00010110","11010101","11100101","00000111","00000000","10110000","11000110","11010000","11000110","11100000",
     "11000110","01000101","00010101","00010000","00010110","11010101","11100101","00000111","00000000","00000101","00000111","00010000","00010110","11010101","11100101","00000111",
     "00000000","00010101","00010111","00001000","00100111","00001000","10000101","00001000","11110110","10010000","00010110","11011000","11100000","11011000","11000101","00010000",
     "11100101","00000111","00000000","11000101","00100111","00000110","11000000","00010111","11000110","00000111","01000000","11011111","01000101","00010111","11100101","00010111",
     "00000111","11000000","00010110","00000111","11000101","01010111","11010111","00010110","11010101","00000111","00010000","11100101","00000111","00000000","00010110","00000111",
     "00100110","00000111","10000101","00000111","11110111","00010110","10010000","11010101","11111000","00100110","00000110","00110110","00000110","10010000","11000000","00000110",
     "11110110","11010110","01000101","00000111","00010000","00010110","11010101","11011111","00010111","00010111","00000111","00000110","00010110","00001000","01011111","00010111",
     "00010110","00000110","00000110","01100110","00000111","01011111","00010101","00010111","00000110","00100111","00000110","00000111","11011111","11000101","00100111","00000110",
     "11000000","00010111","11110110","00000110","01010000","01011111","00000000","11011111","00000111","01110000","00011111","01100000","10011111","00000110","00110000","11011111",
     "00000111","00000000","00011111","00100000","10011111","00001000","01110000","11011111","00000111","01010000","00011111","00000110","01000000","01011111","00000001","10000001",
     "10010001","00100001","00110001","01000001","01100001","01110001","00010001","01010001","00000101","00000101","00000001","00000001","10000001","00000100","00000100","00000100",
     "00000100","00000100","00000100","00000100","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000101","00000110","00000110","00000111",
     "00000111","00000101","11000001","00000100","00001010","01011111","00000001","00100101","10100111","11000001","00000101","00000111","00010111","11110101","00000111","10000001",
     "01110100","00000100","01110100","11000000","00000100","01100101","11010101","11100111","11000001","00100111","11110001","01110111","00000111","01100101","11010101","00100111",
     "11110001","01110111","00000100","10000001","11000001","00000111","00000100","00001010","10011111","00000001","00100101","10100111","11000001","00000101","00000111","00010111",
     "11110101","00000111","10000001","01110100","11000000","00000100","01000111","11010111","11100100","11000001","00100100","10000001","01110100","00000001","00000100","00000100",
     "00001001","01000100","01001111","00000101","00001001","01001001","01001111","00000101","10000100","11000001","10000001","01000001","00000001","11000001","10000001","01000001",
     "00000001","11000001","00000001","00000000","00100100","10000001","01110100","10011111","10100100","01110100","11011111","00000101","01011111","00000001","10010001","00010001",
     "11111111","10000001","00100001","00110001","01000001","01010001","01100001","01110001","10000001","10010001","10100001","10010111","00000101","00010101","10100000","00000101",
     "00000111","00100110","00000110","00000110","00011000","00000101","00000110","00001001","00000101","00000000","00101000","11001110","00000101","00000111","00100111","11011001",
     "11010111","11000111","00011000","00010101","10000011","00000100","01011111","10000000","00100100","00001100","00001100","00000000","00101111","10111110","00000101","00001000",
     "00000111","01000110","00100111","11100110","11010110","10110111","00011110","01000101","01101000","00001110","00000111","10011111","01001100","00001101","00000000","00000000",
     "00000000","00000000","00111111","00010011","00001110","10000000","00000101","01000110","00000101","00000111","00010110","00000110","00000101","00000101","11100111","11100110",
     "10100101","11110101","11000100","00000101","01000110","00000101","00000000","00000111","00010110","00011110","11101110","00001110","00000110","10011111","00000000","00001111",
     "00000101","00001100","00101011","00001100","00001000","00001011","00000011","00000000","00000110","00000111","00100111","00100110","00000111","11100110","11011000","10100111",
     "01001000","00100011","10101000","00001100","00000000","00000000","00000000","00000000","00001110","00000000","11000000","00000101","00010110","00000101","01001000","00000111",
     "10000110","00001000","00000101","00000101","11100111","11100110","10100101","11110101","11010100","00001000","00010110","00000101","00000000","01001000","00000111","10000110",
     "00010011","01001110","10000011","00001111","00000101","00001100","00001100","00000000","00001011","00001111","00000000","00001000","00000101","00001110","00000000","00000000",
     "00000110","00001000","00010111","00100110","11000111","00101000","11110110","11011000","10000111","00010011","01001000","00100101","10000011","00011111","00101110","01001111",
     "10001111","00001100","00000000","00000000","00000000","00000000","00001110","00000000","11000000","00000101","00010110","00000101","01001000","00000111","10000110","00001000",
     "00000101","00000101","11100111","11100110","10100101","11110101","11010100","00001000","00010110","00000101","00000000","01001000","00000111","10000110","00010011","01001110",
     "10000011","10001111","00000101","00000000","00001011","00001100","00000000","00001110","00001110","00001100","00000000","00000000","00000011","00001000","00010110","00101000",
     "11100111","00100011","00100111","01010111","11110111","11110111","11110111","11111000","00001110","10000110","00010101","01001110","00101110","10000101","00010110","00101100",
     "01001100","10000110","00000000","00000000","00000000","00000000","00001010","00000000","11000000","00000101","00010110","00000101","01001000","00000111","10000110","00001000",
     "00000101","00000101","11100111","11100110","10100101","11110101","11010100","00001000","00010110","00000101","00000000","01001000","00000111","10000110","00010011","01001010",
     "10000011","10001111","00000000","00001011","00000000","00000111","00100111","00010110","00110111","11100111","10000110","00010110","00101011","10000110","11000001","10000001",
     "00000101","01000001","00000001","11000001","10000001","01000001","00000001","11000001","10000001","01000001","00000001","00000101","00000001","00000000","00000000","00001111",
     "00000101","00000000","01001111","00000101","00000000","10001111","00000101","00000000","11001111","01011111","00000001","10000001","00010001","00000110","00000101","10000101",
     "11000101","01000101","00000101","10011111","00000100","10000001","11000001","00000001","11001111","00000001","10000001","10010001","00100001","00000101","00000110","00010000",
     "11110101","11000011","01000011","00000000","00001000","00000000","00000111","00010101","11100111","00110111","00000111","10100101","00000101","00010010","01010100","00000101",
     "00000001","00010101","00000011","00000000","00010000","01110100","11111110","00001111","00000000","00000110","00001000","00000111","10111110","00100101","00011000","00011000",
     "11110110","00000111","11100110","11000110","11100110","11000111","00000111","00000111","11110111","11100101","11110111","11110011","10101000","00011111","10001111","10101111",
     "01010011","11110111","11000001","11000111","01000111","10010110","00100110","01110110","11110110","10000001","01000001","00000001","00000000","01100011","11110000","11110000",
     "00100000","11011111","00000101","00000101","10100000","00100101","00010101","00101110","00000000","00000000","00000000","00000000","00111110","00011111","00001110","10000000",
     "00000101","01000111","00000101","00000110","11111000","00000111","00000101","00000101","11010111","11010101","10100101","11100101","10110110","00001000","01000111","00000101",
     "00000000","00000110","11111000","00010011","11011110","01101111","00000000","00000000","00000000","00000101","10100000","00010101","00011110","00100101","00000110","00000000",
     "00101110","11011000","00000101","00000011","00000111","01000110","00100111","11010111","11100110","11111000","00011000","11100101","11000011","00010101","00000000","00000101",
     "10100000","00010101","00000110","11010101","00011000","00000110","00000000","00101000","11010011","00001000","00000111","00100111","11100110","11100111","11110110","00010101",
     "00011000","10110101","00000000","00000101","00010101","00100101","10100101","11010110","00000101","00000110","00000110","00000000","00001000","00000111","00100111","00101000",
     "00010111","11100101","10100101","11110011","01000101","11010110","11000101","00000000","00000101","00010101","00000001","10000001","00000110","01100110","00100101","00000101",
     "01100110","00000000","00000110","00000010","00001000","00001110","00001111","00000000","00000111","00000101","00100111","01100101","00000111","11100110","11001000","11111110",
     "00101110","01001000","11011111","00010011","01101111","01101110","10000010","01110101","11000001","00000001","00000000","00000000","00000101","00010101","00000001","10000001",
     "00000110","01100110","00100101","00000101","01100110","00000000","00000110","00000010","00001000","00001110","00001111","00000000","00001000","00000110","00100110","01101000",
     "11100111","00100111","01010111","11110111","11110111","11110111","11110101","10111000","11001110","00101110","01001000","11011111","00010011","01101111","01101110","10000010",
     "01110101","11000001","00000001","00000000","00000000","11110000","00000101","11000011","11110111","00000111","00000101","00000110","11110110","11100110","10110111","10110111",
     "10110111","10110111","00000111","11010111","00000110","00000000","11000011","00100110","00000000","01010110","11000110","10110111","10110111","10110111","10110111","10110111",
     "10110111","10110111","10110111","10110111","10110111","10110111","10110111","10110111","10110111","10110111","00000000","11110101","10000101","11010101","00000101","11010101",
     "11011111","00100111","00000000","01010110","00000000","00000110","00000010","00000111","11110111","11110110","11000011","11011111","00000001","00000000","00010001","10000001",
     "10010001","00100001","00110001","01000001","01010001","01100001","01110001","10000001","10010001","10100001","10110001","11111111","00000001","00000111","11000111","00100111",
     "00000101","10100001","11110111","11100001","00011111","00010000","00001111","10100001","00100000","01001111","10100001","00110000","10001111","10100001","01000000","11001111",
     "10100001","01010000","00001111","00000101","10100001","00000000","00000111","11111111","00100111","11110111","11110001","11000111","00000111","00010000","11100111","01000001",
     "00000111","00000111","01000001","00010101","01010111","11110111","01100000","11110111","11000001","00000000","00001000","00101000","11111111","10111000","00100111","00000001",
     "00010111","11100000","10110001","00000101","00000001","01000111","11000110","00000101","00010101","00000101","00000101","00000000","10100110","11111111","00000000","10100001",
     "00000110","00000111","00000101","00000110","00000111","01000111","00000111","00000000","00000111","11111111","00100111","11110111","00000001","11000111","01000001","11110001",
     "00011111","10000001","00000111","00010000","11110001","00000000","11111111","00000111","11000100","00100111","10010111","10000001","00000000","00100111","11100111","00010111",
     "11110001","01011111","10000001","00000001","00000001","00001001","00010000","00000100","00011111","01000001","01001111","10100001","11110000","00000100","10011111","01000001",
     "11001111","10100001","00000100","00010100","10001001","10011111","11011111","01011111","00000101","10100000","10100111","10000001","00010111","11100111","11110001","00000000",
     "10000101","01011111","00011111","00000000","11111111","00000100","00100111","11000100","10100111","10011111","01011111","10011111","00000100","00100111","10000111","00000101",
     "11000111","00000101","00000000","11110001","11011111","01000001","00000101","11100111","11011111","01000001","00000101","00000111","11011111","00000101","01000001","00011111",
     "00000000","01010111","00000101","11110101","10100111","00000000","00101001","11110101","00000000","01010111","11110101","00000000","00000000","10000101","01111010","00000000",
     "10011111","10101001","10000001","01001010","00000000","10001100","00000000","00000000","00000110","00000000","00000111","11111111","00100111","11010111","11110001","00000000",
     "01000000","01000001","10110100","00100110","11010111","11011101","11000110","01010110","00011101","00001000","10001100","00000100","00000111","00000100","00001101","00001010",
     "11001101","01001101","01000001","10110100","00100100","10010111","10011101","11000100","00000100","00010110","00000110","01100100","01000110","00000000","00001010","00001101",
     "01000111","01011111","11000100","00010110","11010100","01000001","10110100","00100100","10010111","10011101","11000100","00100110","00000110","10000100","10000110","10000001",
     "00000000","00001101","01000111","11011111","11000100","11000100","00010110","11000100","01000110","00000110","01000001","10110100","00100100","10000111","10001101","10100100",
     "00100110","11000100","01011111","01000001","00000111","00000111","01000001","01100000","11110111","11011111","00000000","00000111","00100111","11111111","11110111","11000111",
     "10000111","11110001","11001111","11000001","10100001","00100111","00000111","00000000","00000111","00100111","11111111","11110111","11110001","01000001","11100111","01000001",
     "11000111","11000111","00000111","11000111","01000001","00001111","11000001","10011111","00000000","00100111","11110101","00000000","11111010","11110101","00000000","01000101",
     "10001010","00000000","00000000","11011111","01001001","10000001","10011010","01011111","00000000","00001001","00001101","10000111","10011111","11000100","00010110","00000110",
     "00000110","11010100","01011111","00000001","11110100","00000000","11011111","01000001","10100100","00000000","10000101","11011111","00000000","00001011","00000101","11011111",
     "00001011","00001011","10011111","00000101","00000000","10000101","00011111","00000100","00001011","00001011","00000100","01011111","00000101","00001011","00001011","01011111",
     "10010000","10100111","10001100","10000001","00000000","10000101","11110101","00000100","00000100","01011111","00000000","00000000","00000101","11000101","00011111","00000000",
     "00000000","01000101","00000101","11011111","00000000","00000000","10000101","00000101","10011111","00000000","00001001","10000101","10011111","11000001","00010111","00000110",
     "10001100","00000110","00000000","00000111","11111111","00100111","11110111","00000000","00000000","11110001","00000000","01000100","01000001","10000111","00100111","11110111",
     "11111001","01100111","00000100","01001001","10011111","00010100","10001100","00000100","00000100","11110100","11000001","00100111","00000110","10001100","00000110","00000000",
     "00000111","11111111","00100111","11110111","00000000","00000000","11110001","00000000","01000100","01000001","10000111","00100111","11110111","11111001","10000111","00000100",
     "00001001","01011111","00010100","10001100","00000100","00000100","11110100","11000001","01000111","00000111","10001100","00000111","00000000","00000111","11111111","00100111",
     "11110111","00000000","00000000","11110001","00000000","01000100","01000001","10000111","00100111","11110111","11111001","10100111","00000100","11001001","00011111","00010100",
     "10001100","00000100","00000100","11110100","00000000","10001100","00000111","11111111","00100111","00000000","00000000","00100111","00000000","00000111","01000100","10000111",
     "00100111","11111001","11111001","01000111","00000100","10001010","00011111","00010100","10001100","00000100","00000100","11110100","00000100","10010000","00000000","00000101",
     "10011111","11100001","00001111","00000001","11000001","00000000","10000001","01000001","00000001","11000001","10000001","01000001","00000001","11000001","10000001","01000001",
     "00000001","11000001","00000001","00000000","01110000","11110001","11011111","00000000","00000110","00100110","00000110","00000001","11000001","00000110","00010000","00000111",
     "11000000","10100110","00000001","11000101","11000001","00000110","00011111","10100110","00000001","11111111","00010110","00000110","00000110","00000011","00000000","00000011",
     "00100011","00010011","00010001","00001000","00000101","00011111","00000000","01000101","10011111","00011111","10100001","00010000","11111001","00010000","00011111","00000000",
     "01000101","01011111","11011111","00000000","10000101","01011111","00010100","11011111","10001100","10000001","00001011","00001011","11110100","11001111","10100100","00000000",
     "00000101","01011111","11011111","01000111","00000111","11011111","00000000","00000000","10000101","10011010","00000000","00000000","10011111","11111001","10000001","00001010",
     "00011111","00000000","00000000","10000101","00101010","00000000","00000000","11011111","01111001","10000001","00001010","01011111","00000000","10000101","00011111","00000000",
     "01110000","00000000","01001001","11110001","01110000","00011010","10011111","00000000","10011111","00000110","00000110","00000101","00000101","00000110","11000101","00000001",
     "11100110","00000000","11110110","10000110","10000000","11111111","00000111","11010111","00000111","11110111","00000000","11110111","00000111","11100101","11110101","11100110",
     "00000111","11100101","00001000","11001000","00001000","00000110","00000011","11001000","10100110","00000111","11110111","10111000","00011000","11110101","00011000","10111000",
     "00000111","10111000","11001000","00000011","00000011","11001000","11100110","00001000","01101000","11011000","00001000","11110111","00011000","11100111","11011000","00000111",
     "00000101","11100101","00000000","00000000","00000110","00010000","11000111","00000001","11101000","00000000","11111000","10001000","10000000","11111111","00000111","11010111",
     "00000111","11110110","00000000","11010111","00000111","00001000","00010101","00001000","00001110","00010000","00000011","11100111","11100111","11010101","00000111","11110111",
     "11010111","00010111","11110101","00010111","11010111","00000111","11010111","11100111","00000011","00000011","11100111","11010111","00000111","01100111","11010111","11111000",
     "11110111","00010111","11100111","11010111","00000110","00000101","11100101","00000000","11010101","00000001","11110110","00000000","11110110","10000110","10000000","11111111",
     "10000111","11100111","00000111","00000000","00000111","11101110","00001110","10110110","11000101","00010101","00000000","00000000","00000000","00000000","00000000","11110000",
     "11010111","10000110","10000000","00011111","11110000","00001000","00010111","10001000","10000000","00011111","11110000","00000110","11000111","10000110","10000000","10011111",
     "11111000","11010101","00001000","11100110","11110101","11010101","11100110","00001000","00001110","11110101","00000111","11100110","11001110","00000110","10110110","11110110",
     "00010110","11111110","00010110","11110110","11101110","00010110","11110110","11100110","00000111","00000111","11100110","11001110","00000110","11110111","10100111","00010111",
     "11110110","00010111","10100111","11100110","00010111","00001110","10100111","11000101","10011111","11100110","11000110","11010111","11100101","00000110","11100011","00000110",
     "00001110","11000101","11100101","00000111","00001000","11000110","11100011","11111110","00000011","00010011","10111000","11011000","11110111","11011000","10111000","11100111",
     "11011000","10111000","11101000","00001000","00001000","11101000","11101110","00001000","00001000","01100101","11010101","11110111","11010101","01100101","11100111","11010101",
     "00000111","00000001","11100111","11111111","11100111","00000111","11100110","00000110","11100110","01100101","11000110","00001110","11101000","11100110","11011000","11001000",
     "11100110","11100110","00000110","11001000","11000101","11000101","00000111","00000000","00000000","00000001","11110111","11100110","00000110","11101110","11000101","11010110",
     "11010101","11110111","00000000","00000000","00000110","00000000","01011111","00000110","00000000","00011111","00001000","00000000","01011111","00000000","00010000","00000000",
     "00000110","00000000","01011111","00001000","00011111","00000111","11011111","00000111","01011111","00000110","00011111","11100101","00011000","00011111","11100101","00010111",
     "10011111","10100101","00110111","11000101","00000111","00110000","11000111","00110101","00000101","00000111","11001000","00000110","11110111","11000111","00000101","00000111",
     "00000110","01000111","01000110","00000111","11000111","11110110","11100111","11000111","01000111","11110111","11110101","00010111","00000000","00000101","00010101","00000101",
     "00010111","00010101","11110111","00010111","00000000","00000101","00010111","00110111","11010111","00010101","00000111","00000101","00010111","00110111","11010111","00010101",
     "00000111","01011111","00000101","01000101","10000101","11000101","00000101","01000101","10000101","11000101","01000101","11010111","11000101","01010111","11110111","11100111",
     "11010111","11000111","01100111","00000111","01000111","11010111","11110111","10011111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
  signal ram_symbol3 : ram_type := (
     "10000000","00001011","00000000","00000000","00000000","00000000","00000000","00000000","11111110","11111110","11111110","11111110","11111110","11111110","11111110","11111110",
     "11111100","11111100","11111101","11111101","11111101","11111101","11111101","11111101","11111100","00010101","00000011","00000011","00000011","00000011","00000010","00000010",
     "00000010","00000010","00000001","00000001","00000001","00000001","00000000","00000000","00000000","00000000","00000100","00110000","00000000","01011110","00000000","01001000",
     "00000000","11011110","10000011","00000000","00000000","00000000","11111111","00000000","10100100","11111111","00000000","10100011","00000000","00000000","00000000","00000000",
     "00000000","00000000","11111110","00000000","00000000","10001000","00110000","00000000","10000000","00110000","00100100","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","00110011","00110111","01100010","01100110","01101010","01101110","01110010","01110110","01111010",
     "00000000","00110011","00110111","01000010","01000110","01001010","01001110","01010010","01010110","01011010","00000000","01001100","00000000","01010010","01110110","01110010",
     "01110011","00100000","01101110","00100000","00100101","01111010","00000000","01010010","01110110","01111000","01110100","00100000","01100101","01101011","01110101","01100101",
     "01101001","00101001","01101000","01101101","01110100","00100000","01100101","01101101","00101110","00000000","01001111","00110010","01101100","01100101","01110100","01101110",
     "01100101","01101111","00100000","01110111","01100101","01110100","01110010","01110010","00001010","00000000","01110010","01101001","00001010","00000000","01110000","01101111",
     "01101110","01110010","01110000","01101101","01110010","01101111","01101111","01100001","00001010","00000000","01110110","01100100","01101111","01110101","01100001","01100101",
     "01110011","01110010","01110010","01110010","00000000","01100110","00100000","01100101","01101001","01110010","01110000","01101101","01110010","01101111","01101111","01100001",
     "00001010","00000000","01110000","01101111","01101110","01110010","01110000","01101101","01110010","01101111","01101111","01100001","00001010","00000000","01110110","01100100",
     "01101111","01110101","01100001","01100101","01110011","01110010","01110010","01110010","00000000","01011101","01001111","01101100","00100000","00100000","00110000","00101101",
     "01101111","00100000","00110000","00110100","00000000","01011101","01001111","01101101","01101001","01110010","01111000","01111000","01110011","01101100","01100101","00100101",
     "00001010","00000000","01011101","01001111","01110011","01100101","01100011","00100101","00100000","01101000","01100100","00100000","00110000","00000000","01100101","01101011",
     "01111010","00100000","00100101","00000000","01100001","01101001","00100000","00100000","00100101","00000000","01100001","01101001","00101000","01110011","00100101","00000000",
     "01110010","01101111","01010011","00100000","00100101","00000000","01001111","01001101","00100000","01100011","00100000","00100000","01101100","01110100","00100000","01110011",
     "01110010","01110110","01100100","01110011","00100001","00000000","01110010","01101111","00100000","00100000","00100101","00000000","00111000","00110000","00000000","01110000",
     "01110010","01110010","01101110","00100101","00000000","01100100","01110101","00100000","00100000","01100101","01100101","00000000","01110000","01110010","01100001","00100000",
     "00100101","00000000","01000011","00000000","01101111","01101100","01110100","00100000","00100101","00000000","01100100","00100000","00100000","00100000","00110000","00110100",
     "00000000","01011101","01101100","00100000","00100000","00100000","00110000","00000000","01011101","01101101","01101001","00100000","00100000","00110000","00000000","01011101",
     "01110011","01100101","00100000","00100000","00110000","00000000","01011101","01100110","01101100","00100000","00100000","00110000","00000000","01110010","00100000","01110010",
     "01101111","01100001","01100001","00101110","01100101","01000001","00101110","01100110","01110010","01100001","01110010","01110010","01100111","01101100","00001010","00000000",
     "01101111","01100100","01100011","00001010","00000000","01101110","01110110","01100100","00100000","01110010","01101111","01101111","01101000","00100000","01100100","01101100",
     "00101100","01100101","00100000","01110000","00100000","01101000","01110011","01110011","00100000","01101110","00100000","01110100","01101101","00000000","01110100","00000000",
     "01110000","00000000","01100011","00000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000",
     "10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","10000000","00110011","01000110","00000000","01010100","01110001","00000000","00101110",
     "01111010","00000000","00110000","01011110","00000000","00110000","00110011","00000000","00110010","00110010","00000000","01100101","00110010","00000000","00110110","00110010",
     "00000000","00110101","00110000","00000000","00110011","00110000","00000000","00110000","00110000","00000000","00110110","00110000","00000000","00110010","00000000","00110100",
     "00000000","00110100","00000000","00110010","00000000","00000010","00000011","00000100","00000100","00000101","00000101","00000101","00000101","00000110","00000110","00000110",
     "00000110","00000110","00000110","00000110","00000110","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111",
     "00000111","00000111","00000111","00000111","00000111","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000","00001000",
     "00001000","00001000","00001000","00001000","00001000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000100","10000000","01010100","00000000","00000000","00000000","00000000","10000000","11101011","00000000","10000010","00000000","10000010",
     "00000000","10000000","11101001","00000000","10000010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00001111","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00001111","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00001111","00000001","00000000","00000001","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00001111","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000001","00000000","00001111","00000001","00000000","00000001","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00001111","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00001111","00000001","00000000","00000001",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00001111",
     "00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000",
     "00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","11111111",
     "00000000","00000000","00000001","00000001","00000000","00000000","00000000","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00000000","11110110",
     "00001000","00001001","00001000","00001000","00001001","00001001","00001001","00001001","00000111","00000111","00000111","00000111","00000111","00000100","00000000","00000000",
     "00011110","10000000","01111000","00000001","00011100","00000000","00000001","00000011","00011010","00000000","00000010","00011100","00011100","00000000","00100000","00000000",
     "00000000","00000000","11111111","00000010","00000000","00000001","00100000","11111111","00000000","01000000","00011010","00000011","00000000","00000000","00000000","00000000",
     "00000001","00000000","00000000","00000000","01000001","11111111","00000010","00011111","00000000","00000000","00000010","00000000","01110010","00000000","00000001","11111111",
     "11111111","00000000","00000000","00000000","00000000","00000000","00011010","00000001","00010110","00000010","00011011","11111111","01000001","00000001","00000000","11111111",
     "00000000","00000000","00000000","01000001","01101100","00000001","11111111","00000001","01000001","00000000","00000000","00000011","01101010","00000001","00000001","00000000",
     "00000000","00000000","00000000","01000000","00000001","11111110","00000000","11111111","11111110","00000001","00000011","11111111","01000001","00000000","00000000","00000000",
     "00000000","00000010","01100100","00000000","00001001","00001001","00000000","00001001","00001001","00001000","00001000","00001000","00001000","00000111","00000111","00000111",
     "00000111","00000110","00001010","00000000","11111111","00000000","00000000","00000010","00000010","00000000","11100100","10000000","01110101","11100001","00000000","11100101",
     "01000000","11111111","00000010","11100100","00000000","00000001","00000000","00000000","00000011","00000000","00000001","00000000","00000000","00000000","00000000","00000011",
     "11111110","11111101","11100011","11111111","00000010","11011111","00000011","00000000","00000111","00000000","00000000","11100111","11111111","11011111","00000011","00000000",
     "00000000","11100110","00000000","11111111","11101000","11111111","00000000","00000000","11100010","00000000","00000010","11110000","00000000","00000001","00001111","11111110",
     "00000000","00000000","11110000","00000000","00000001","00001111","11111110","00000000","00000000","11111100","11100111","00010101","00010110","00010110","00010110","00010111",
     "00010101","00010101","00010101","00010101","00010101","00010101","00010101","00010011","00010110","00010110","00010110","00011000","00011000","00011001","00011001","00000000",
     "00010111","00000001","00100110","00000011","10000000","10000000","10000000","00000000","00000000","01010101","01011001","01110101","10000000","00000010","00001010","00000000",
     "00000000","00000000","00000000","11111110","00000000","00000011","01000000","00000000","00000000","11110000","00000000","01000001","00000110","00000000","00000001","00001111",
     "11111110","00000000","00000000","00000000","00000000","11111100","00010110","00010110","00010110","00010110","00010101","00010101","00010101","00010101","00010100","00010100",
     "00010100","00010100","00010011","00011001","00000000","00000000","00000001","00001111","11111110","00000001","11111000","00000000","00000001","00000000","11111110","00001111",
     "00000000","00000010","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","11111110","00001111","11111100","11111101","00001111","00000000",
     "00001100","00000010","11111111","00001110","00000010","11111111","00001000","00001101","00000100","00000100","11111011","00001111","00000011","00101010","00000000","00000001",
     "00000000","00000000","00000001","00000000","11111001","00000000","00000000","11111000","00000010","00000000","11110111","00000000","00000000","11110110","00000000","00000011",
     "00000000","11111011","00001111","00100110","10000000","00000000","01100111","00000000","00000000","00000000","00000000","00000000","00000000","11111101","00001111","00100110",
     "00000010","00101000","00000000","00000000","11110100","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111101","11111101","00001111",
     "11111100","11110000","00000000","00000000","00000000","00000000","11101110","01000000","00000001","11101110","00000000","00000100","00000001","00000000","00000000","00000000",
     "00000000","10011111","00000000","00000000","00000000","11011010","11011011","00000000","00000000","11111101","00000000","00000000","00000000","01101000","00000000","00001000",
     "00001000","00000000","00000000","01000000","00000000","00000000","00000000","11111110","00000001","01000000","01100100","00001010","00000000","00000000","00000000","00000000",
     "11111111","00000000","00000000","00000000","00000000","00000000","00000000","00000110","00000000","00000000","00000110","11111111","00000000","00000000","00000000","00000000",
     "00000000","00000000","11111110","11111110","11111111","00000000","00000000","00000000","00000010","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","01000000","00000000","00000000","00000010","00001110","00000000","00000000","11001000","11001001","00000000",
     "11111111","01010100","00000000","00000001","00000000","11101010","00000000","00000000","11101001","00000000","00000001","11111111","01010010","00000000","00000000","00000000",
     "00000000","00000000","01110110","00000000","00000010","00000000","00000111","00000000","00000000","11000000","11000010","00000000","00000000","00000010","00000000","01001010",
     "00000000","00000000","01001000","00000000","00000000","00000011","11000000","00000000","11000011","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","11111101","11111101","00001111","11111100","00000000","11001100","00000000","00000000","00000000","11111111","01000001","00000000","00000000","11001010","00000110",
     "00000000","00000000","00000000","11011011","00111111","00000110","00000000","00000100","00000000","01011000","10000000","01111000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000000",
     "00000000","00000001","00000001","00000001","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000011","00000000","00000000","00000000","00000000","00000010","00000010","00000010","00000000","00000000","00000001","00000001","00000001",
     "00000011","00000010","00000011","00000011","00000000","00000010","00000000","00000001","11111111","00000010","01000010","00000001","01000010","11111110","00000000","00000010",
     "00000000","00000000","01101000","00000001","00000001","00000000","01011110","00000000","00000000","00000000","00000000","00000000","10100000","10100001","00000110","00000000",
     "00000000","01000010","00000000","11101010","00000000","00000001","11000001","00000000","00000000","00000000","00110000","00000110","01001000","00000110","00000010","00000000",
     "00000000","00000000","00000000","00000010","00000011","00000000","00000000","00000000","00000000","00000000","00000011","00000000","00000000","00000000","00010011","00000000",
     "11101110","00010011","00000000","00000000","00000010","11101111","00101100","00000110","00111100","00000110","00000000","00010011","00000000","00000000","00000011","00000011",
     "00000011","00000000","00000000","11101110","00000001","00000000","00000011","11101111","00000000","00000000","00010011","00000000","00000000","11101110","00010011","00000000",
     "00000000","00000010","11101110","00000000","00100110","00000110","00110010","00000110","00000000","00010011","00000000","00000000","00000011","00000011","00000011","00000000",
     "00000000","11101110","00000001","00000000","00000011","11101111","00000000","00000000","00010011","00000000","00000000","11101110","00000000","00010011","00000000","00000010",
     "11101110","00000000","00100010","00000110","00110000","00000110","00000000","00010011","00000000","00000000","00000010","00000010","00000011","00000000","00000000","11101110",
     "00000000","00000000","00000011","11101110","00000000","00000000","00010011","00000000","00000000","11101110","00000001","11111111","00000010","00110110","01000000","00000000",
     "00000000","00000010","00000000","01000100","00000000","00000001","01000000","00000001","11111111","00000000","00000000","00000001","00000000","00111001","00000000","00000000",
     "00000000","00000010","00000010","00000000","00000000","01000001","00000001","11111110","00000000","11111110","00000000","00000000","11111000","11111001","00000000","00000000",
     "00000000","00000000","00000000","00000000","10011011","00000000","00000100","00000000","11011000","00000000","00000000","00000000","00000001","00000000","00000000","00000000",
     "11110010","11110100","00000000","00000000","10101011","00100100","00000000","00000000","00000010","00000000","00110110","11111111","10101100","01111010","10011000","11111111",
     "00100100","01000000","00000000","00000000","00000010","00000000","00110011","00000000","00000001","01000000","00000001","10011000","00000011","00000000","00000000","00010011",
     "00000000","00000000","00000010","11101111","00000000","11010100","00010011","00000000","00000011","11101110","00000000","00010011","00000000","00000000","00000010","11101110",
     "00000000","11011000","00010011","00000000","00000011","11101110","00000000","00010011","00000000","00000000","00000010","11101110","00000000","11011100","00010011","00000000",
     "00000011","00000000","11101110","11100001","11111111","00000000","00000000","00000001","00000001","00000000","00000000","00011101","00000000","00000001","00000001","10111110",
     "00000010","00000001","00000001","00000000","01000000","00000000","11111110","00000000","11111110","10111100","00000011","00000000","11011110","00000000","10111110","00000000",
     "11010000","00000000","00000011","00010011","00000000","00000000","00000000","00000000","00000011","11101110","11001111","00000000","11000110","00000000","00000011","00010011",
     "00000000","00000000","00000000","00000000","00000011","11101110","11000100","00000000","11010010","00000000","00000010","00010011","00000000","00000000","00000000","00000000",
     "00000010","11101110","11010000","00000000","00000010","00000000","00000011","00000000","00000000","00000000","00000000","00000000","00000011","00000000","10110111","00000000",
     "00000000","00000000","10110110","00000001","11011110","00000000","10000011","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11001010","11001101",
     "00000000","11110110","00000000","00000000","11111111","00000000","11111110","11111110","11111110","11111111","00000000","00000000","11001011","11111110","00000001","00000000",
     "00000000","00000000","00000001","00000000","01000000","00000000","00000111","00000100","00000000","01000000","00000000","00000000","00000000","00000000","00000000","00000011",
     "00000100","00000000","00001000","00000001","00000001","00000000","00000000","00000111","11110000","11100011","00000000","00000010","00001000","00000000","00000001","00000001",
     "00000000","00000001","00000001","00000000","00000010","00000000","00000010","00000000","00000000","00000010","00000000","00000000","00000001","00000001","00001111","01001111",
     "00000011","00000001","01000001","00000000","00000010","00000011","11111000","00000000","00000010","00111100","00000011","00000001","01000001","11111110","00000011","00000010",
     "11110101","11111110","00000000","00000001","00000001","00000000","00000000","00000001","00000000","00000000","00000000","01000000","00000000","00000111","00000100","01000000",
     "00000000","00000000","00000000","00000000","00000000","00000011","00001100","00000000","00010100","00000001","00000001","00000000","00000000","00000111","11110000","11010010",
     "00000000","00000010","00001000","00000000","00000000","01000000","00000000","00000111","00000100","01000000","00000000","00000000","00000000","00000000","00000011","00001010",
     "00000000","00010000","00000001","00000001","00000000","00000000","00000111","11110000","11001011","00000000","00000010","00001000","00000000","00000001","00000001","01000001",
     "00000001","00000001","00000000","00000000","00000010","00000000","00000010","00000000","00000000","00000010","00000000","00000000","00000001","00000001","00001111","00110111",
     "00000011","00000001","01000001","00000000","00000010","00000011","11110001","00000010","00000000","00000000","00000010","00000000","00000000","00000001","00000001","00001111",
     "00110011","00000011","00000001","01000001","00000000","00000010","00000011","11110011","00000000","00000010","00100000","00000011","00000001","01000001","11111000","00000011",
     "00000010","11101010","00000000","00000010","00011101","00000011","00000001","01000001","11111010","00000011","00000010","11101110","00000000","00000000","00000000","01000000",
     "00000000","00000000","00000001","00000001","00000000","11110000","00000000","00000000","00000000","00000001","00000001","00000000","11110000","00000000","00000000","00000000",
     "00000000","01000000","00000000","00000000","00000000","00000000","00000000","00000000","11111010","00000011","00000100","00000100","00000100","00000101","00000101","00000101",
     "00000101","00000101","00000011","00000011","00000011","00000011","00000000","00000000","00000000","00000010","00111001","00000000","00000000","00000000","00000000","00000000",
     "00000000","00001111","00000000","00101010","01011110","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000",
     "11111110","00000000","00000000","00000000","00000000","00000000","00000000","11111110","00101000","00000000","00000000","00000001","00000000","00000001","00000000","00000000",
     "01000000","00000000","00000000","00000001","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000001",
     "01000001","00000000","00000000","00000001","01000001","11110010","00000000","01000001","00000000","00000001","00000001","00000000","00101000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00010010","00000000","00000000","00000000","00000000","00000000","11111110",
     "00000000","00000010","00000000","00000001","00000000","10010001","00000000","00000000","11111110","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111110","00000000","00000000","00000000",
     "00000000","00000110","00001010","00001010","00000000","00000000","00000000","00000001","00000001","00000000","11110000","00000001","00000000","00000000","00000000","00000001",
     "00000001","11110000","00000000","00000001","00000000","00000000","01000001","00000110","00000000","00000000","11111111","00000010","00000000","00000000","11111000","00000100",
     "00000100","00000000","11111111","00000000","11111110","00000000","00000000","11111101","00000000","00000001","00000000","11101100","00000000","11111110","00000000","11101100",
     "11101110","00000000","11111111","00000000","11111001","11110000","00000000","00000111","00000000","00101000","00000000","00000000","00000000","00000000","11101110","00110100",
     "00000000","00000000","00000000","00000000","11010111","00000000","00000001","00000000","11010110","00000000","11111110","11010101","00000000","00000000","00000001","00000000",
     "00000001","00000000","00000000","00000001","00000001","11011001","00000000","00101110","00000000","00000001","00000000","11110100","00000000","00000000","11111110","00000101",
     "00000101","00000101","00000101","00000100","00000100","00000100","00000100","00000011","00000011","00000011","00000011","00000010","00000110","00000000","00000000","00000000",
     "11010110","00011010","00000000","00000000","00000010","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","11111110","00000000","00001110","00010000","00010000","00000000","00000000","00000000","00001000","00000111","00000100","01000000",
     "00000000","00000000","00000000","00000000","00000011","00011010","00011001","00000001","00000001","00000000","00000000","11101011","00000111","11110000","00000001","00000010",
     "00001000","00000001","00000000","00001000","00000111","00000100","01000000","00000000","00000000","00000000","00000000","00000011","00001110","00001011","00000001","00000001",
     "00000000","00000000","11100101","00000111","11110000","00000001","00000010","00001000","00000001","01000000","00000100","00000000","00000000","11111111","00000010","00000000",
     "00000000","11110000","00000010","00000010","00000000","11111111","00000000","11111110","00000000","00000000","11111101","00000000","11111111","00000000","11111100","00000000",
     "11101010","00000001","00000000","00000000","10111110","00000000","00000000","00000000","11100110","00000000","00000000","00000001","00000000","00111011","00000011","00000001",
     "01000001","00000100","00000011","00000010","11110011","00000010","00000000","00000000","00000010","00000000","00000000","00000001","00000001","00001111","01001000","00000011",
     "00000001","01000001","00000000","00000010","00000011","11101111","00000001","00000000","00110100","00000011","00000001","01000001","00000100","00000011","00000010","11100110",
     "00000010","00000000","00000000","00000010","00000000","00000000","00000001","00000001","00001111","01000001","00000011","00000001","01000001","00000000","00000010","00000011",
     "11100010","00000001","11010011","00000000","00000000","00000001","00000010","00000000","11111111","00001000","00000001","00000000","11111111","00000000","00000001","00000001",
     "00000000","00000000","00000000","00000001","00000001","00000000","00100011","00000000","00000000","00100011","00000000","00000001","00000000","11111111","11111111","00000000",
     "00000000","00000000","00000110","00000001","11111111","00000001","00000000","11111111","00000000","00000101","00000000","00000101","00000001","00000001","00000000","00000000",
     "00000111","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111011","00000000",
     "00000010","00000000","00000010","00000000","00000000","11111111","00000000","00010010","00000000","00000000","00000000","00000000","11111110","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000000","00000000","00000110","00001000","00001000",
     "00000000","00000000","00000000","00000001","00000001","00000000","11110000","00000000","00000001","00000000","00000000","00000001","00000001","11110000","00000000","00000001",
     "00000001","00000000","01000000","00000100","00000000","00000000","11111111","00000010","00000001","00000000","11111000","00000010","00000010","00000000","11111111","00000000",
     "11111110","00000000","00000000","11111101","00000000","11111111","00000000","11111100","11110010","00000000","00000100","00000000","11110000","00000000","00000000","00000001",
     "00000001","00000000","00000000","01110000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","11101010","11101100","00000000","00000000","00000000",
     "00000000","00000000","11100000","00000000","00000000","11011111","00000000","00000000","00000100","00000000","00000000","00000100","00000001","00000000","00000000","00000001",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000010","00000010","00000000","00000000","00000000","00000101","00000000","00000000","00000000","00000000","11111110","00000000","11111110",
     "00000000","00000000","00000000","00000000","00000010","00000000","00000000","00000000","00000000","11111110","11111101","00000000","00000000","00000000","00000010","00000000",
     "00000000","00000000","00000000","00000000","00000000","11111110","00000000","00010100","11111101","00000001","00000001","00000001","00000001","00000001","00000010","00000010",
     "00000010","00000011","00000001","00000001","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","11111111","00000000","00000010","00000100","00000100","00000000","00000000","00000000","00000000","00000100","00000000","00000000",
     "11111111","00000010","00000000","00000000","11111100","00000010","00000010","00000000","11111111","00000000","11111110","00000000","00000000","11111101","00000000","11111111",
     "00000000","11111100","00000000","11110110","00000000","00000001","00000000","11110100","00000000","00000000","00000010","00000010","00000000","00000010","00000010","00000001",
     "00000001","00000001","00000001","00000000","00000000","00000000","00000000","00000011","00000000","00000000","00000000","00000000","00000000","00000000","10000000","00000000",
     "00000000","11101010","11101010","11110000","00000100","00000000","00000100","00000000","00100100","00000000","11111111","00000100","00000000","00000100","00000000","11110000",
     "00000100","10000000","11101010","11101010","00000000","10000000","10000000","11101010","11101011","11101010","11101011","01000000","00000000","01000000","01000000","00000000",
     "11111111","00000110","00000000","00000000","01000001","00000000","00000001","00000000","11111111","00000000","00000000","10000000","00000110","01111011","00000000","11000010",
     "10000000","00000000","01111101","11000001","00000000","00000000","00000000","00000000","00000001","00000000","00000000","10000000","10000010","10111111","00000000","11111111",
     "00000000","00000000","00000000","00000001","00000001","00000010","00000010","00000000","00000000","00000100","00000000","00000000","10110011","00000011","11100110","00000010",
     "11111111","00000000","10110001","00000011","11100100","00000010","00000010","00000000","11111100","00000000","00000000","00000000","00000000","00000000","00000001","00000000",
     "00000010","00000000","11111100","00000000","11111001","00000000","00000010","11110000","00000000","00000001","00001111","11111110","00000000","00000000","00000000","11111110",
     "00000000","00000000","00000010","11110000","00000000","00000001","00001111","11111110","00000000","00000000","00000000","11111110","11110000","00000000","00000001","00001111",
     "11111110","00000000","00000000","00000000","11111111","00000000","00000000","00010100","00000000","00000001","00000001","00000000","11111111","00000001","10000000","10000000",
     "00000000","00000000","00000001","00000000","11001010","11001001","00000000","00000010","00000000","00001010","00000000","00000001","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000001","00000001","00000001","00001010","00000000","00000000","00000001","00000000","00000000","00000001","00000000","00000001","00000000","00000001",
     "00000010","00000000","00000001","00000000","00000001","00000000","00000001","00000001","00000000","00000000","00000000","00000001","00000000","11111111","00000001","00000000",
     "00000001","00000000","00000000","11110100","00000000","00000000","00000000","00000001","00000000","00000000","00000001","00000000","00000000","11110110","00000001","00000010",
     "00000001","11110100","00000010","01000001","00000000","00000001","01100111","00000001","00000011","00000001","11110010","11111110","00000000","00000000","01000001","00000000",
     "00000001","01100101","00000000","00000000","00101110","00000010","00000000","00101011","00000000","11111101","00001111","00000000","00000000","00001010","00000001","00000000",
     "00010110","00000000","00010101","11111101","00000010","00000000","00000010","00001111","00000011","00001100","00000000","00000000","00000000","00010010","00101010","00000000",
     "11111101","00001111","11111101","00000001","00000000","00000000","00000000","00101000","00000010","00000000","00100010","00000100","00000000","00000010","11111101","00001101",
     "00001111","00001111","00011010","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000010","00000100","00000010","00000100","00000010",
     "00011000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000001","00000000","00011100","00000000","00011011","00000000","11111101","00001111","00000000","00000000","00000010","00000010","00010100","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000010","00000000","11101010","00000000","00000000","11111000","00000001","00000000","00000000","00000000",
     "00010010","00000010","00000000","00010011","00000000","11111101","00001111","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00001110",
     "00000000","00001111","00000001","11111101","00001111","00000000","00000000","00000000","11111100","00000000","00001010","00000000","00001011","00000000","00000010","11111101",
     "00001111","00000000","00000000","00000000","00000000","00000000","00000000","11101101","00000000","00000000","00000000","00000110","00001011","00000000","11111100","00000000",
     "00000000","00000000","00000100","00000100","00000000","11100010","00000001","00000000","00000010","00000000","00000011","00000000","11011111","00000000","00000000","00000000",
     "00000010","00000000","11111110","00000000","00000000","11100110","00000000","11100101","00000000","00000000","11100101","00000000","11100100","00000000","00000000","11100011",
     "00000000","00000000","11100011","00000000","11100010","00000000","00000000","11100001","00000000","00000000","11100001","00000000","00000000","11100000","11111000","00000110",
     "00000110","00000111","00000111","00000111","00000111","00000101","00000110","00000111","00000000","00000000","00000011","00000010","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000010","00000010","00000010","00000010","00000000","00000000","00000000","00000000",
     "00000000","00010100","00000000","00000000","00000000","11000011","00000101","00000000","00000000","00000000","11111100","00000000","00000000","11111100","11111100","00000000",
     "00000001","00000000","00010011","00000010","00000000","00000001","00000010","00000000","00000000","00000001","00000000","00000001","00000000","00000001","11111110","00000001",
     "00000000","11111111","00000000","00000000","00000000","00000010","00000000","00000000","10111010","00000101","00000000","00000000","00000000","11111100","00000000","00000000",
     "11111100","11111100","00000000","00000011","00000010","00000000","00000001","00000110","00000000","00000000","00000001","00000000","11111111","00000001","00000000","00000000",
     "00000000","00000000","10011101","00000000","00000000","00000000","10011100","00000000","11111100","00000111","00000111","00000111","00000111","00000110","00000110","00000110",
     "00000110","00000101","00001000","00000000","00000001","00000000","11110111","11111001","00000000","11101111","11111000","11110010","11111000","11111101","00000010","00000010",
     "11111111","00000010","00000011","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000001","00000000","01001000","00000000","01000000","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "11111110","11111110","00000000","01000001","00000000","00000000","11111101","01000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000010","11111110","11111110","00000000","00000001","01000000","00000001","00000000","11111100","00000001","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000001","00000000","00000001","00000001","00000000","01000001","00000000","00000011","00000000","00000001","00000001","00000000","00000000",
     "00000000","00000000","11111100","00000001","00000000","01000001","00000000","00000000","11111101","00000000","01000001","00000001","00000000","11111001","00000000","11001111",
     "00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000011","00000000","00000000","11111110",
     "00000000","00000001","11111101","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000001","00000000","01000001","00000000","00000000",
     "00000100","00000000","00000001","00000001","00000000","00000000","00000000","00000000","11111100","00000001","00000000","01000001","00000000","00000000","00000000","11111100",
     "00000000","00000001","11111000","11000010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000011","00000001","00000000","00000000","11111110","00000000","00000000","00000000","11111010","00000000","00000001","00000001",
     "11111010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000001","00000000","01000001","00000000","00000000","00000100","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","11111100","00000001","00000000","01000001","00000000","00000000","00000000","11111100","00000000","00000001",
     "11111000","10110010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000010","00000001","01000000","01000000","00000000","00000111","00000010","00000000","00000001","11111100","00000000","00000000","00000000","11111010","00000000","00000001",
     "00000001","11111000","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000001","00000000","01000001","00000000","00000000","00000100","00000000",
     "00000001","00000001","00000000","00000000","00000000","00000000","11111100","00000001","00000000","01000001","00000000","00000000","00000000","11111100","00000000","00000001",
     "11111000","10100010","00000000","00000000","00000000","00000000","00000000","00000000","01000001","11111110","11111110","00000000","00000001","11111100","00000010","00000010",
     "00000001","00000010","00000010","00000001","00000001","00000001","00000001","00000000","00000000","00000000","00000000","01000001","00000011","00000000","00000000","10011011",
     "00000000","00000000","10011010","00000000","00000000","10011001","00000000","00000000","10011000","11111001","11111111","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","10101110","00000000","00000000","00000000","00000001","10010100","11111111","00000000","00000000","00000001","00000000","00000000","00000000",
     "11111111","11111111","00000000","00000000","00000000","00001110","00000000","00000000","00000010","00000000","11111111","00000010","00000000","00000000","00000000","00001000",
     "00000000","00000000","00000000","00000000","00000000","01000000","11111111","00000000","00000000","00000011","00000001","00000001","00000000","00000000","00000000","00000000",
     "01000001","00000001","00000000","00000001","01000000","00000000","00000001","00000001","00000000","11111110","00001111","00000000","11111010","00000000","00000000","11111010",
     "00000000","11111111","00000000","11111111","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000001","00000000","00000000","11111111","11111111",
     "00000000","11110011","00000000","00001000","01000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000001","00000000","00000001",
     "00000001","00000000","01000001","00000000","00000010","00000000","00000001","00000001","00000000","00000000","00000000","00000000","11111100","00000001","00000000","01000001",
     "00000000","00000000","11111100","00000000","01000001","11111010","00000000","00000000","00000000","00000100","01000000","00000000","00000000","00000000","00000001","00000000",
     "00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000010","11111110","11111110","00000000","00000001","01000001","11111101","00000000","00000100",
     "01000000","00000000","00000001","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111110","11111110","00000000",
     "01000001","11111100","00000000","00000100","00000000","00000000","00000000","00000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000011","00000000","00000000","11111110","00000000","00000001","11111101","00000000","00001000","00000000","11111111","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000011","00000000","00000000","11111110",
     "00000000","00000000","11111101","00000000","00000000","00000000","00000000","11111010","00000000","00000001","00000000","00000000","00001010","00000000","11111111","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000010","01000000","01000000","00000000","00000111","00000010","00000000","00000000","11111100","00000000","00000000","11111011","00000000","00000000","00000000","00000000",
     "11111000","00000000","00000001","00000000","00000000","00000000","00000000","00000010","00000000","00001010","00001000","11111111","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000001","11111110","00000000","00000000","01000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00001111","00000000","00000000","00000001","00000000",
     "11110110","00000000","00000000","00000000","00000000","11111010","00000000","11111111","01000000","00000000","11110110","11110011","10000001","00000000","01111110","01111110",
     "01111110","01111111","01111101","01111101","01111101","01111101","01111101","01111101","01111101","01111101","01111011","11111111","11111000","10000011","01111101","00000000",
     "00000000","00000000","00000000","00000101","11011001","00000000","10101111","00000000","00000000","10101110","00000000","00000000","10101101","00000010","00000000","10101100",
     "00000010","00000000","10101100","01111100","00000010","00000000","10000011","11111111","00000000","00000000","00000000","01111110","00111000","00000000","00000010","00000000",
     "01111111","00000000","00000000","00110100","01000001","01111110","00000110","01111110","00000011","00000000","10000011","00000000","11111111","00000000","00000000","00000110",
     "00000000","00000000","00000000","01111111","00000100","00000000","00000000","00000000","00000000","00000001","00000001","01111101","00000010","11111111","00000000","00000010",
     "01110000","01110100","01110010","00110000","00110100","00000000","00000010","00000000","10000011","11111111","00000000","00000000","00000011","01111110","00000011","00000000",
     "11011101","00000011","00001010","00000000","00000010","00000000","11111111","10000011","01111110","00000000","00000000","00000011","00000000","00000000","00000000","00000000",
     "00000010","10110111","00000011","00000100","00000100","00000100","00000000","00000000","11111100","00000101","10101111","00000100","11111111","00000000","11111010","00000101",
     "10101101","00000100","01101110","00000000","11111100","10110110","10110111","10111010","11111000","00000000","00000010","00000011","00000000","00000010","00000010","10000000",
     "10000110","11111110","10101111","00000000","11111111","10000011","00000000","01111110","00000000","10111101","10110001","10110010","10000011","00000000","00000000","00000000",
     "01111110","00000000","00000000","00000000","10011101","00000000","00000000","01111110","10011100","00000000","00000000","01111111","10011011","00000000","00000011","10011011",
     "00000000","10110000","00000000","01101000","00100000","00000000","10100000","01101010","00000000","10011111","00100110","10000000","00000000","10010000","11111101","00000000",
     "11110010","11100011","00000001","01110001","10000000","11101001","00000000","00000000","01101010","00000000","10000011","11111111","00000000","00000000","00000000","00000000",
     "00000100","00000000","00000001","00000000","00000000","00000000","10000010","00000001","00000000","00000001","11101001","00000001","00000001","00000001","00000001","01000001",
     "00011100","00000000","00000000","00000001","00000000","00000000","00000000","10000000","10000010","00000000","00000010","10000010","00000011","10000000","00000000","00000000",
     "10010110","11100110","10000010","00000000","10000010","00000000","00000001","00000000","00000000","00000000","10000000","00000000","00000010","10000010","00000011","00000000",
     "10000000","00000000","10011001","11100001","10000010","10000000","00000000","10000010","00000000","11110010","00000000","00000001","00000000","00000000","00000000","10000010",
     "00001111","10000010","11110001","00000000","01111111","11001000","00000000","00000110","01111110","11000111","00000000","10000011","00000000","11111111","00000000","01111110",
     "01111111","00000000","10111000","00000011","00000100","00000000","11001010","00000000","10000011","00000000","11111111","00000000","00000000","00000000","01111110","00000011",
     "01111110","01111111","00000001","00000000","00000100","11100101","00000011","11000111","00000000","10001111","01001100","00000000","11101010","00000100","10000000","10001101",
     "01100000","00000000","00000000","11010001","01011010","00000001","10100111","11011111","10000000","00000000","00000000","10011100","11001111","10000010","00000000","00000001",
     "00000001","10000010","11100001","00000000","11111111","10000000","10011001","00000011","00000000","10000000","10011111","11001011","10000000","00000000","10100001","11001010",
     "00000000","00000000","10000011","00000000","10000000","10100010","11001001","00000001","00000000","00000000","00000001","10000001","00110110","00000000","00000000","10000000",
     "00000000","00110100","11101001","00000011","10000000","10101001","00000010","00000001","01000001","11000100","10000000","10000000","10101011","10101011","11000011","10000000",
     "10000000","10101101","10101111","11000001","10000000","10000000","10110000","10110001","11000000","10000000","00000000","10110010","10111111","00000011","00000000","00000110",
     "11101001","00000110","00000000","10000011","11111111","00000000","00000000","00000000","10000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","10000010","00000000","10110100","10111001","00000000","11101001","00000001","00000001","11111100","00000011","00000000","00000110","11101001","00101000","00000000",
     "10000011","11111111","00000000","00000000","00000000","10000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10000010","00000000",
     "10110110","10110010","00000000","11101001","00000001","00000001","11111100","00000011","00000000","00000110","11101001","00001100","00000000","10000011","11111111","00000000",
     "00000000","00000000","10000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","10000010","00000000","10110111","10101011","00000000",
     "11101001","00000001","00000001","11111100","00000000","11101001","10000011","11111111","00000000","00000000","10000000","00000001","00000000","00000010","00000000","00000000",
     "00000000","00000000","00000000","10000010","00000000","10111001","10100101","00000000","11101001","00000001","00000001","11111100","00010000","00001110","10000000","11000000",
     "10100010","00000101","11100010","00001000","01111110","00000000","01111110","01111110","01111110","01111101","01111101","01111101","01111101","01111100","01111100","01111100",
     "01111100","01111011","01111111","00000000","00000000","00000010","10000011","00000000","10000011","00000000","00000001","00000110","00000000","01111111","00000000","10001100",
     "00000001","00000010","00000110","00000000","00000010","10001010","10111101","00000010","00000110","11111111","00000000","00000001","00000001","00000001","00000000","10000011",
     "00000000","00000001","00000001","01111111","10000110","11111011","10000000","11000001","10010100","11110010","00000100","00000000","10010010","00000000","10001110","10000000",
     "10111011","10010010","11101111","10000000","10100101","10010001","00000000","11001010","11101001","00000011","00000000","00000000","00000010","11001000","00000010","10000000",
     "10100100","10001110","11000110","00000000","11100100","11101001","10000000","00000000","10001010","00011001","00000000","00000000","10001011","10011011","00000001","00110100",
     "10011001","10000000","00000000","10000111","11100101","00000000","00000000","10001000","11100100","00000001","01001011","10010110","10000000","10010011","10000111","00000000",
     "01110100","00000000","11011000","00000000","01110100","00111100","10010011","00000000","10110111","00000000","00000000","00000000","00000000","00011010","00001100","00000000",
     "00100010","00000001","01000000","00000001","00000001","11111111","10000000","00000000","00000000","00000000","00000010","01000000","00000000","00000000","00000000","00000000",
     "00000001","00000000","00000001","00000010","00000001","00000001","00000001","00000010","00000010","00000001","00000000","00000000","00000001","11111111","00000001","00111110",
     "00000000","01000000","00000010","00000001","00000001","00000010","00000010","00000001","00000000","00000000","00000001","11111111","00000001","11111111","00000000","00000000",
     "00000001","00000000","00000000","00000000","00000000","00000000","00000010","00000000","00010010","00000001","00110100","00000001","00000001","11111111","01110010","00000000",
     "00000000","00000000","00000010","01000000","00010010","00000001","01000001","00000001","00000001","00000000","00000001","00000011","00000011","00000011","00000001","00000000",
     "00000000","00000001","11111111","00000001","00110010","00000000","01000000","00000011","00000001","00000001","00000011","00000011","00000001","00000000","00000001","00000000",
     "11111111","00000001","11111111","00000001","00000000","00000001","00000000","00000000","00000100","00000000","00000100","00000001","00100110","00000001","00000001","11111111",
     "01100101","00000000","00000000","00000010","00000001","01000000","00010000","00100100","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00001111",
     "00100100","00000000","00000000","11111011","00001111","00000000","11101101","00000000","00000000","11101101","00001111","00000000","11011110","00000000","00000000","11011101",
     "00000000","00000000","00000001","00000011","00000000","00000000","00000000","00000001","00000001","00000000","00000001","00000011","00000011","00000001","00000000","00000000",
     "00000001","11111111","00011101","00011100","11111111","00000001","01000000","00000011","00000001","00000001","00000011","00000010","00000001","00000000","00000000","00000001",
     "11111111","00011001","00011000","11111111","00000001","00000001","01000000","00000000","11100100","00000000","00000001","00000000","00000000","00000001","00000011","00000001",
     "00000001","00000001","00000000","00000001","00000001","00000001","00000011","00000010","00000001","00000001","00000000","00000000","11111111","00010010","00010010","11111111",
     "00000000","01000000","00000011","00000001","00000001","00000011","00000010","00000001","00000001","00000000","00000000","11111111","00001100","00001100","11111111","00000000",
     "00000001","00000000","00000000","11111111","00000000","00000001","00000000","00000001","00000010","01000000","00000010","00000001","00000010","00000000","00000000","00000010",
     "00000000","00000001","00000001","00000000","00000010","00000000","00000000","00000000","00000000","00000000","11111111","00000000","00000001","00000000","00000001","00000001",
     "11111100","11111111","00000000","00000000","00000001","00000001","11011010","00000001","00000001","10111111","00000001","00000001","11001100","00000000","00000000","00000000",
     "00000000","00000000","11010111","00000000","11110011","00000000","11100111","00000000","11101110","00000000","11100011","11111111","00000001","11000001","11111111","00000001",
     "11001101","00000000","00000000","00000000","00000110","00000000","00000100","00000000","00000000","00000110","11111111","11111110","00001000","00000010","00000000","00000000",
     "00000000","00000000","00000000","11111111","11111110","11111111","01000000","11111111","00000000","00000000","00000000","00000001","00000000","00000000","11111111","00000000",
     "00000000","00000000","11111110","11111111","00000000","00000000","00000000","00000000","11111110","00000000","11111000","00000000","00000000","00000000","11111110","00000000",
     "11111100","11110110","00000000","00000000","00000000","00000000","00000001","00000001","00000001","00000001","00000010","00000000","11111111","00000000","00000001","00000001",
     "00000001","00000001","00000000","00000001","00000010","11111110","11111010","11110001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000");
  signal zz_1 : std_logic_vector(7 downto 0);
  signal zz_2 : std_logic_vector(7 downto 0);
  signal zz_3 : std_logic_vector(7 downto 0);
  signal zz_4 : std_logic_vector(7 downto 0);
begin
  zz_Axi4Incr_result_1 <= pkg_extract(Axi4Incr_base,11,1);
  zz_Axi4Incr_result_2 <= pkg_extract(Axi4Incr_baseIncr,0,0);
  zz_Axi4Incr_result_3 <= pkg_extract(Axi4Incr_base,11,2);
  zz_Axi4Incr_result_4 <= pkg_extract(Axi4Incr_baseIncr,1,0);
  zz_Axi4Incr_result_5 <= pkg_extract(Axi4Incr_base,11,3);
  zz_Axi4Incr_result_6 <= pkg_extract(Axi4Incr_baseIncr,2,0);
  zz_Axi4Incr_result_7 <= pkg_extract(Axi4Incr_base,11,4);
  zz_Axi4Incr_result_8 <= pkg_extract(Axi4Incr_baseIncr,3,0);
  zz_Axi4Incr_result_9 <= pkg_extract(Axi4Incr_base,11,5);
  zz_Axi4Incr_result_10 <= pkg_extract(Axi4Incr_baseIncr,4,0);
  zz_Axi4Incr_result_11 <= pkg_extract(Axi4Incr_base,11,6);
  zz_Axi4Incr_result_12 <= pkg_extract(Axi4Incr_baseIncr,5,0);
  process (zz_1, zz_2, zz_3, zz_4)
  begin
    zz_ram_port0 <= zz_4 & zz_3 & zz_2 & zz_1;
  end process;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if stage0_fire = '1' then
        zz_1 <= ram_symbol0(to_integer(zz_io_axi_r_payload_data));
        zz_2 <= ram_symbol1(to_integer(zz_io_axi_r_payload_data));
        zz_3 <= ram_symbol2(to_integer(zz_io_axi_r_payload_data));
        zz_4 <= ram_symbol3(to_integer(zz_io_axi_r_payload_data));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_axi_w_payload_strb(0) = '1' and stage0_fire = '1' and stage0_payload_fragment_write = '1' then
        ram_symbol0(to_integer(zz_io_axi_r_payload_data)) <= zz_io_axi_r_payload_data_1(7 downto 0);
      end if;
      if io_axi_w_payload_strb(1) = '1' and stage0_fire = '1' and stage0_payload_fragment_write = '1' then
        ram_symbol1(to_integer(zz_io_axi_r_payload_data)) <= zz_io_axi_r_payload_data_1(15 downto 8);
      end if;
      if io_axi_w_payload_strb(2) = '1' and stage0_fire = '1' and stage0_payload_fragment_write = '1' then
        ram_symbol2(to_integer(zz_io_axi_r_payload_data)) <= zz_io_axi_r_payload_data_1(23 downto 16);
      end if;
      if io_axi_w_payload_strb(3) = '1' and stage0_fire = '1' and stage0_payload_fragment_write = '1' then
        ram_symbol3(to_integer(zz_io_axi_r_payload_data)) <= zz_io_axi_r_payload_data_1(31 downto 24);
      end if;
    end if;
  end process;

  process(Axi4Incr_wrapCase,zz_Axi4Incr_result_1,zz_Axi4Incr_result_2,zz_Axi4Incr_result_3,zz_Axi4Incr_result_4,zz_Axi4Incr_result_5,zz_Axi4Incr_result_6,zz_Axi4Incr_result_7,zz_Axi4Incr_result_8,zz_Axi4Incr_result_9,zz_Axi4Incr_result_10,zz_Axi4Incr_result_11,zz_Axi4Incr_result_12)
  begin
    case Axi4Incr_wrapCase is
      when "000" =>
        zz_Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(zz_Axi4Incr_result_1),std_logic_vector(zz_Axi4Incr_result_2)));
      when "001" =>
        zz_Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(zz_Axi4Incr_result_3),std_logic_vector(zz_Axi4Incr_result_4)));
      when "010" =>
        zz_Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(zz_Axi4Incr_result_5),std_logic_vector(zz_Axi4Incr_result_6)));
      when "011" =>
        zz_Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(zz_Axi4Incr_result_7),std_logic_vector(zz_Axi4Incr_result_8)));
      when "100" =>
        zz_Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(zz_Axi4Incr_result_9),std_logic_vector(zz_Axi4Incr_result_10)));
      when others =>
        zz_Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(zz_Axi4Incr_result_11),std_logic_vector(zz_Axi4Incr_result_12)));
    end case;
  end process;

  unburstify_buffer_last <= pkg_toStdLogic(unburstify_buffer_beat = pkg_unsigned("00000001"));
  Axi4Incr_validSize <= pkg_extract(unburstify_buffer_transaction_size,1,0);
  Axi4Incr_highCat <= pkg_extract(unburstify_buffer_transaction_addr,14,12);
  Axi4Incr_sizeValue <= unsigned(pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_unsigned("10") = Axi4Incr_validSize)),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_unsigned("01") = Axi4Incr_validSize)),pkg_toStdLogicVector(pkg_toStdLogic(pkg_unsigned("00") = Axi4Incr_validSize)))));
  Axi4Incr_alignMask <= pkg_resize(unsigned(pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_unsigned("01") < Axi4Incr_validSize)),pkg_toStdLogicVector(pkg_toStdLogic(pkg_unsigned("00") < Axi4Incr_validSize)))),12);
  Axi4Incr_base <= (pkg_resize(pkg_extract(unburstify_buffer_transaction_addr,11,0),12) and pkg_not(Axi4Incr_alignMask));
  Axi4Incr_baseIncr <= (Axi4Incr_base + pkg_resize(Axi4Incr_sizeValue,12));
  process(unburstify_buffer_len)
  begin
    if (pkg_toStdLogic((std_logic_vector(unburstify_buffer_len) and pkg_stdLogicVector("00001000")) = pkg_stdLogicVector("00001000")) = '1') then
        zz_Axi4Incr_wrapCase <= pkg_unsigned("11");
    elsif (pkg_toStdLogic((std_logic_vector(unburstify_buffer_len) and pkg_stdLogicVector("00001100")) = pkg_stdLogicVector("00000100")) = '1') then
        zz_Axi4Incr_wrapCase <= pkg_unsigned("10");
    elsif (pkg_toStdLogic((std_logic_vector(unburstify_buffer_len) and pkg_stdLogicVector("00001110")) = pkg_stdLogicVector("00000010")) = '1') then
        zz_Axi4Incr_wrapCase <= pkg_unsigned("01");
    else
        zz_Axi4Incr_wrapCase <= pkg_unsigned("00");
    end if;
  end process;

  Axi4Incr_wrapCase <= (pkg_resize(Axi4Incr_validSize,3) + pkg_resize(zz_Axi4Incr_wrapCase,3));
  process(unburstify_buffer_transaction_burst,unburstify_buffer_transaction_addr,Axi4Incr_highCat,zz_Axi4Incr_result,Axi4Incr_baseIncr)
  begin
    case unburstify_buffer_transaction_burst is
      when "00" =>
        Axi4Incr_result <= unburstify_buffer_transaction_addr;
      when "10" =>
        Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(Axi4Incr_highCat),std_logic_vector(zz_Axi4Incr_result)));
      when others =>
        Axi4Incr_result <= unsigned(pkg_cat(std_logic_vector(Axi4Incr_highCat),std_logic_vector(Axi4Incr_baseIncr)));
    end case;
  end process;

  process(unburstify_buffer_valid,unburstify_result_ready)
  begin
    io_axi_arw_ready <= pkg_toStdLogic(false);
    if unburstify_buffer_valid = '0' then
      io_axi_arw_ready <= unburstify_result_ready;
    end if;
  end process;

  process(unburstify_buffer_valid,io_axi_arw_valid)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_valid <= pkg_toStdLogic(true);
    else
      unburstify_result_valid <= io_axi_arw_valid;
    end if;
  end process;

  process(unburstify_buffer_valid,unburstify_buffer_last,when_Axi4Channel_l181)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_payload_last <= unburstify_buffer_last;
    else
      if when_Axi4Channel_l181 = '1' then
        unburstify_result_payload_last <= pkg_toStdLogic(true);
      else
        unburstify_result_payload_last <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

  process(unburstify_buffer_valid,unburstify_buffer_transaction_id,io_axi_arw_payload_id)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_payload_fragment_id <= unburstify_buffer_transaction_id;
    else
      unburstify_result_payload_fragment_id <= io_axi_arw_payload_id;
    end if;
  end process;

  process(unburstify_buffer_valid,unburstify_buffer_transaction_size,io_axi_arw_payload_size)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_payload_fragment_size <= unburstify_buffer_transaction_size;
    else
      unburstify_result_payload_fragment_size <= io_axi_arw_payload_size;
    end if;
  end process;

  process(unburstify_buffer_valid,unburstify_buffer_transaction_burst,io_axi_arw_payload_burst)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_payload_fragment_burst <= unburstify_buffer_transaction_burst;
    else
      unburstify_result_payload_fragment_burst <= io_axi_arw_payload_burst;
    end if;
  end process;

  process(unburstify_buffer_valid,unburstify_buffer_transaction_write,io_axi_arw_payload_write)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_payload_fragment_write <= unburstify_buffer_transaction_write;
    else
      unburstify_result_payload_fragment_write <= io_axi_arw_payload_write;
    end if;
  end process;

  process(unburstify_buffer_valid,Axi4Incr_result,io_axi_arw_payload_addr)
  begin
    if unburstify_buffer_valid = '1' then
      unburstify_result_payload_fragment_addr <= Axi4Incr_result;
    else
      unburstify_result_payload_fragment_addr <= io_axi_arw_payload_addr;
    end if;
  end process;

  when_Axi4Channel_l181 <= pkg_toStdLogic(io_axi_arw_payload_len = pkg_unsigned("00000000"));
  zz_unburstify_result_ready <= (not (unburstify_result_payload_fragment_write and (not io_axi_w_valid)));
  stage0_valid <= (unburstify_result_valid and zz_unburstify_result_ready);
  unburstify_result_ready <= (stage0_ready and zz_unburstify_result_ready);
  stage0_payload_last <= unburstify_result_payload_last;
  stage0_payload_fragment_addr <= unburstify_result_payload_fragment_addr;
  stage0_payload_fragment_id <= unburstify_result_payload_fragment_id;
  stage0_payload_fragment_size <= unburstify_result_payload_fragment_size;
  stage0_payload_fragment_burst <= unburstify_result_payload_fragment_burst;
  stage0_payload_fragment_write <= unburstify_result_payload_fragment_write;
  zz_io_axi_r_payload_data <= pkg_extract(stage0_payload_fragment_addr,14,2);
  stage0_fire <= (stage0_valid and stage0_ready);
  zz_io_axi_r_payload_data_1 <= io_axi_w_payload_data;
  io_axi_r_payload_data <= zz_ram_port0;
  io_axi_w_ready <= ((unburstify_result_valid and unburstify_result_payload_fragment_write) and stage0_ready);
  process(stage1_ready,when_Stream_l342)
  begin
    stage0_ready <= stage1_ready;
    if when_Stream_l342 = '1' then
      stage0_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Stream_l342 <= (not stage1_valid);
  stage1_valid <= stage0_rValid;
  stage1_payload_last <= stage0_rData_last;
  stage1_payload_fragment_addr <= stage0_rData_fragment_addr;
  stage1_payload_fragment_id <= stage0_rData_fragment_id;
  stage1_payload_fragment_size <= stage0_rData_fragment_size;
  stage1_payload_fragment_burst <= stage0_rData_fragment_burst;
  stage1_payload_fragment_write <= stage0_rData_fragment_write;
  stage1_ready <= ((io_axi_r_ready and (not stage1_payload_fragment_write)) or ((io_axi_b_ready or (not stage1_payload_last)) and stage1_payload_fragment_write));
  io_axi_r_valid <= (stage1_valid and (not stage1_payload_fragment_write));
  io_axi_r_payload_id <= stage1_payload_fragment_id;
  io_axi_r_payload_last <= stage1_payload_last;
  io_axi_r_payload_resp <= pkg_stdLogicVector("00");
  io_axi_b_valid <= ((stage1_valid and stage1_payload_fragment_write) and stage1_payload_last);
  io_axi_b_payload_resp <= pkg_stdLogicVector("00");
  io_axi_b_payload_id <= stage1_payload_fragment_id;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      unburstify_buffer_valid <= pkg_toStdLogic(false);
      stage0_rValid <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if unburstify_result_ready = '1' then
        if unburstify_buffer_last = '1' then
          unburstify_buffer_valid <= pkg_toStdLogic(false);
        end if;
      end if;
      if unburstify_buffer_valid = '0' then
        if when_Axi4Channel_l181 = '0' then
          if unburstify_result_ready = '1' then
            unburstify_buffer_valid <= io_axi_arw_valid;
          end if;
        end if;
      end if;
      if stage0_ready = '1' then
        stage0_rValid <= stage0_valid;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if unburstify_result_ready = '1' then
        unburstify_buffer_beat <= (unburstify_buffer_beat - pkg_unsigned("00000001"));
        unburstify_buffer_transaction_addr(11 downto 0) <= pkg_extract(Axi4Incr_result,11,0);
      end if;
      if unburstify_buffer_valid = '0' then
        if when_Axi4Channel_l181 = '0' then
          if unburstify_result_ready = '1' then
            unburstify_buffer_transaction_addr <= io_axi_arw_payload_addr;
            unburstify_buffer_transaction_id <= io_axi_arw_payload_id;
            unburstify_buffer_transaction_size <= io_axi_arw_payload_size;
            unburstify_buffer_transaction_burst <= io_axi_arw_payload_burst;
            unburstify_buffer_transaction_write <= io_axi_arw_payload_write;
            unburstify_buffer_beat <= io_axi_arw_payload_len;
            unburstify_buffer_len <= io_axi_arw_payload_len;
          end if;
        end if;
      end if;
      if stage0_ready = '1' then
        stage0_rData_last <= stage0_payload_last;
        stage0_rData_fragment_addr <= stage0_payload_fragment_addr;
        stage0_rData_fragment_id <= stage0_payload_fragment_id;
        stage0_rData_fragment_size <= stage0_payload_fragment_size;
        stage0_rData_fragment_burst <= stage0_payload_fragment_burst;
        stage0_rData_fragment_write <= stage0_payload_fragment_write;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4SharedToApb3Bridge is
  port(
    io_axi_arw_valid : in std_logic;
    io_axi_arw_ready : out std_logic;
    io_axi_arw_payload_addr : in unsigned(19 downto 0);
    io_axi_arw_payload_id : in unsigned(3 downto 0);
    io_axi_arw_payload_len : in unsigned(7 downto 0);
    io_axi_arw_payload_size : in unsigned(2 downto 0);
    io_axi_arw_payload_burst : in std_logic_vector(1 downto 0);
    io_axi_arw_payload_write : in std_logic;
    io_axi_w_valid : in std_logic;
    io_axi_w_ready : out std_logic;
    io_axi_w_payload_data : in std_logic_vector(31 downto 0);
    io_axi_w_payload_strb : in std_logic_vector(3 downto 0);
    io_axi_w_payload_last : in std_logic;
    io_axi_b_valid : out std_logic;
    io_axi_b_ready : in std_logic;
    io_axi_b_payload_id : out unsigned(3 downto 0);
    io_axi_b_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_valid : out std_logic;
    io_axi_r_ready : in std_logic;
    io_axi_r_payload_data : out std_logic_vector(31 downto 0);
    io_axi_r_payload_id : out unsigned(3 downto 0);
    io_axi_r_payload_resp : out std_logic_vector(1 downto 0);
    io_axi_r_payload_last : out std_logic;
    io_apb_PADDR : out unsigned(19 downto 0);
    io_apb_PSEL : out std_logic_vector(0 downto 0);
    io_apb_PENABLE : out std_logic;
    io_apb_PREADY : in std_logic;
    io_apb_PWRITE : out std_logic;
    io_apb_PWDATA : out std_logic_vector(31 downto 0);
    io_apb_PRDATA : in std_logic_vector(31 downto 0);
    io_apb_PSLVERROR : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4SharedToApb3Bridge;

architecture arch of Axi4SharedToApb3Bridge is

  signal phase : Axi4ToApb3BridgePhase;
  signal write : std_logic;
  signal readedData : std_logic_vector(31 downto 0);
  signal id : unsigned(3 downto 0);
  signal when_Axi4SharedToApb3Bridge_l91 : std_logic;
begin
  process(phase,io_apb_PREADY)
  begin
    io_axi_arw_ready <= pkg_toStdLogic(false);
    case phase is
      when pkg_enum.SETUP =>
      when pkg_enum.ACCESS_1 =>
        if io_apb_PREADY = '1' then
          io_axi_arw_ready <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  process(phase,io_apb_PREADY,write)
  begin
    io_axi_w_ready <= pkg_toStdLogic(false);
    case phase is
      when pkg_enum.SETUP =>
      when pkg_enum.ACCESS_1 =>
        if io_apb_PREADY = '1' then
          io_axi_w_ready <= write;
        end if;
      when others =>
    end case;
  end process;

  process(phase,write)
  begin
    io_axi_b_valid <= pkg_toStdLogic(false);
    case phase is
      when pkg_enum.SETUP =>
      when pkg_enum.ACCESS_1 =>
      when others =>
        if write = '1' then
          io_axi_b_valid <= pkg_toStdLogic(true);
        end if;
    end case;
  end process;

  process(phase,write)
  begin
    io_axi_r_valid <= pkg_toStdLogic(false);
    case phase is
      when pkg_enum.SETUP =>
      when pkg_enum.ACCESS_1 =>
      when others =>
        if write = '0' then
          io_axi_r_valid <= pkg_toStdLogic(true);
        end if;
    end case;
  end process;

  process(phase,when_Axi4SharedToApb3Bridge_l91)
  begin
    io_apb_PSEL(0) <= pkg_toStdLogic(false);
    case phase is
      when pkg_enum.SETUP =>
        if when_Axi4SharedToApb3Bridge_l91 = '1' then
          io_apb_PSEL(0) <= pkg_toStdLogic(true);
        end if;
      when pkg_enum.ACCESS_1 =>
        io_apb_PSEL(0) <= pkg_toStdLogic(true);
      when others =>
    end case;
  end process;

  process(phase)
  begin
    io_apb_PENABLE <= pkg_toStdLogic(false);
    case phase is
      when pkg_enum.SETUP =>
      when pkg_enum.ACCESS_1 =>
        io_apb_PENABLE <= pkg_toStdLogic(true);
      when others =>
    end case;
  end process;

  when_Axi4SharedToApb3Bridge_l91 <= (io_axi_arw_valid and ((not io_axi_arw_payload_write) or io_axi_w_valid));
  io_apb_PADDR <= io_axi_arw_payload_addr;
  io_apb_PWDATA <= io_axi_w_payload_data;
  io_apb_PWRITE <= io_axi_arw_payload_write;
  io_axi_r_payload_resp <= pkg_cat(pkg_toStdLogicVector(io_apb_PSLVERROR),pkg_stdLogicVector("0"));
  io_axi_b_payload_resp <= pkg_cat(pkg_toStdLogicVector(io_apb_PSLVERROR),pkg_stdLogicVector("0"));
  io_axi_r_payload_id <= id;
  io_axi_b_payload_id <= id;
  io_axi_r_payload_data <= readedData;
  io_axi_r_payload_last <= pkg_toStdLogic(true);
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      phase <= pkg_enum.SETUP;
    elsif rising_edge(io_mainClk) then
      case phase is
        when pkg_enum.SETUP =>
          if when_Axi4SharedToApb3Bridge_l91 = '1' then
            phase <= pkg_enum.ACCESS_1;
          end if;
        when pkg_enum.ACCESS_1 =>
          if io_apb_PREADY = '1' then
            phase <= pkg_enum.RESPONSE;
          end if;
        when others =>
          if write = '1' then
            if io_axi_b_ready = '1' then
              phase <= pkg_enum.SETUP;
            end if;
          else
            if io_axi_r_ready = '1' then
              phase <= pkg_enum.SETUP;
            end if;
          end if;
      end case;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      case phase is
        when pkg_enum.SETUP =>
          write <= io_axi_arw_payload_write;
          id <= io_axi_arw_payload_id;
        when pkg_enum.ACCESS_1 =>
          if io_apb_PREADY = '1' then
            readedData <= io_apb_PRDATA;
          end if;
        when others =>
      end case;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Apb3Gpio is
  port(
    io_apb_PADDR : in unsigned(3 downto 0);
    io_apb_PSEL : in std_logic_vector(0 downto 0);
    io_apb_PENABLE : in std_logic;
    io_apb_PREADY : out std_logic;
    io_apb_PWRITE : in std_logic;
    io_apb_PWDATA : in std_logic_vector(31 downto 0);
    io_apb_PRDATA : out std_logic_vector(31 downto 0);
    io_apb_PSLVERROR : out std_logic;
    io_gpio_read : in std_logic_vector(31 downto 0);
    io_gpio_write : out std_logic_vector(31 downto 0);
    io_gpio_writeEnable : out std_logic_vector(31 downto 0);
    io_value : out std_logic_vector(31 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Apb3Gpio;

architecture arch of Apb3Gpio is
  signal io_apb_PREADY_read_buffer : std_logic;
  signal io_value_read_buffer : std_logic_vector(31 downto 0);
  signal io_gpio_read_buffercc_io_dataOut : std_logic_vector(31 downto 0);

  signal ctrl_askWrite : std_logic;
  signal ctrl_askRead : std_logic;
  signal ctrl_doWrite : std_logic;
  signal ctrl_doRead : std_logic;
  signal io_gpio_write_driver : std_logic_vector(31 downto 0);
  signal io_gpio_writeEnable_driver : std_logic_vector(31 downto 0);
begin
  io_apb_PREADY <= io_apb_PREADY_read_buffer;
  io_value <= io_value_read_buffer;
  io_gpio_read_buffercc : entity work.BufferCC_2
    port map ( 
      io_dataIn => io_gpio_read,
      io_dataOut => io_gpio_read_buffercc_io_dataOut,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  io_value_read_buffer <= io_gpio_read_buffercc_io_dataOut;
  io_apb_PREADY_read_buffer <= pkg_toStdLogic(true);
  process(io_apb_PADDR,io_value_read_buffer,io_gpio_write_driver,io_gpio_writeEnable_driver)
  begin
    io_apb_PRDATA <= pkg_stdLogicVector("00000000000000000000000000000000");
    case io_apb_PADDR is
      when "0000" =>
        io_apb_PRDATA(31 downto 0) <= io_value_read_buffer;
      when "0100" =>
        io_apb_PRDATA(31 downto 0) <= io_gpio_write_driver;
      when "1000" =>
        io_apb_PRDATA(31 downto 0) <= io_gpio_writeEnable_driver;
      when others =>
    end case;
  end process;

  io_apb_PSLVERROR <= pkg_toStdLogic(false);
  ctrl_askWrite <= ((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PWRITE);
  ctrl_askRead <= ((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and (not io_apb_PWRITE));
  ctrl_doWrite <= (((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PREADY_read_buffer) and io_apb_PWRITE);
  ctrl_doRead <= (((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PREADY_read_buffer) and (not io_apb_PWRITE));
  io_gpio_write <= io_gpio_write_driver;
  io_gpio_writeEnable <= io_gpio_writeEnable_driver;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      io_gpio_writeEnable_driver <= pkg_stdLogicVector("00000000000000000000000000000000");
    elsif rising_edge(io_mainClk) then
      case io_apb_PADDR is
        when "1000" =>
          if ctrl_doWrite = '1' then
            io_gpio_writeEnable_driver <= pkg_extract(io_apb_PWDATA,31,0);
          end if;
        when others =>
      end case;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      case io_apb_PADDR is
        when "0100" =>
          if ctrl_doWrite = '1' then
            io_gpio_write_driver <= pkg_extract(io_apb_PWDATA,31,0);
          end if;
        when others =>
      end case;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Apb3UartCtrl is
  port(
    io_apb_PADDR : in unsigned(4 downto 0);
    io_apb_PSEL : in std_logic_vector(0 downto 0);
    io_apb_PENABLE : in std_logic;
    io_apb_PREADY : out std_logic;
    io_apb_PWRITE : in std_logic;
    io_apb_PWDATA : in std_logic_vector(31 downto 0);
    io_apb_PRDATA : out std_logic_vector(31 downto 0);
    io_uart_txd : out std_logic;
    io_uart_rxd : in std_logic;
    io_interrupt : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Apb3UartCtrl;

architecture arch of Apb3UartCtrl is
  signal uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready : std_logic;
  signal io_apb_PREADY_read_buffer : std_logic;
  signal uartCtrl_1_io_write_ready : std_logic;
  signal uartCtrl_1_io_read_valid : std_logic;
  signal uartCtrl_1_io_read_payload : std_logic_vector(7 downto 0);
  signal uartCtrl_1_io_uart_txd : std_logic;
  signal uartCtrl_1_io_readError : std_logic;
  signal uartCtrl_1_io_readBreak : std_logic;
  signal bridge_write_streamUnbuffered_queueWithOccupancy_io_push_ready : std_logic;
  signal bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid : std_logic;
  signal bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_payload : std_logic_vector(7 downto 0);
  signal bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy : unsigned(4 downto 0);
  signal bridge_write_streamUnbuffered_queueWithOccupancy_io_availability : unsigned(4 downto 0);
  signal uartCtrl_1_io_read_queueWithOccupancy_io_push_ready : std_logic;
  signal uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid : std_logic;
  signal uartCtrl_1_io_read_queueWithOccupancy_io_pop_payload : std_logic_vector(7 downto 0);
  signal uartCtrl_1_io_read_queueWithOccupancy_io_occupancy : unsigned(4 downto 0);
  signal uartCtrl_1_io_read_queueWithOccupancy_io_availability : unsigned(4 downto 0);

  signal busCtrl_askWrite : std_logic;
  signal busCtrl_askRead : std_logic;
  signal busCtrl_doWrite : std_logic;
  signal busCtrl_doRead : std_logic;
  signal bridge_uartConfigReg_frame_dataLength : unsigned(2 downto 0);
  signal bridge_uartConfigReg_frame_stop : UartStopType_seq_type;
  signal bridge_uartConfigReg_frame_parity : UartParityType_seq_type;
  signal bridge_uartConfigReg_clockDivider : unsigned(19 downto 0);
  signal zz_bridge_write_streamUnbuffered_valid : std_logic;
  signal bridge_write_streamUnbuffered_valid : std_logic;
  signal bridge_write_streamUnbuffered_ready : std_logic;
  signal bridge_write_streamUnbuffered_payload : std_logic_vector(7 downto 0);
  signal bridge_read_streamBreaked_valid : std_logic;
  signal bridge_read_streamBreaked_ready : std_logic;
  signal bridge_read_streamBreaked_payload : std_logic_vector(7 downto 0);
  signal bridge_interruptCtrl_writeIntEnable : std_logic;
  signal bridge_interruptCtrl_readIntEnable : std_logic;
  signal bridge_interruptCtrl_readInt : std_logic;
  signal bridge_interruptCtrl_writeInt : std_logic;
  signal bridge_interruptCtrl_interrupt : std_logic;
  signal bridge_misc_readError : std_logic;
  signal when_BusSlaveFactory_l335 : std_logic;
  signal when_BusSlaveFactory_l337 : std_logic;
  signal bridge_misc_readOverflowError : std_logic;
  signal when_BusSlaveFactory_l335_1 : std_logic;
  signal when_BusSlaveFactory_l337_1 : std_logic;
  signal uartCtrl_1_io_read_isStall : std_logic;
  signal bridge_misc_breakDetected : std_logic;
  signal uartCtrl_1_io_readBreak_regNext : std_logic;
  signal when_UartCtrl_l155 : std_logic;
  signal when_BusSlaveFactory_l335_2 : std_logic;
  signal when_BusSlaveFactory_l337_2 : std_logic;
  signal bridge_misc_doBreak : std_logic;
  signal when_BusSlaveFactory_l366 : std_logic;
  signal when_BusSlaveFactory_l368 : std_logic;
  signal when_BusSlaveFactory_l335_3 : std_logic;
  signal when_BusSlaveFactory_l337_3 : std_logic;
  function zz_bridge_uartConfigReg_clockDivider return unsigned is
    variable bridge_uartConfigReg_clockDivider : unsigned(19 downto 0);
  begin
    bridge_uartConfigReg_clockDivider := pkg_unsigned("00000000000000000000");
    bridge_uartConfigReg_clockDivider := pkg_unsigned("00000000000010101100");
    return bridge_uartConfigReg_clockDivider;
  end function;
begin
  io_apb_PREADY <= io_apb_PREADY_read_buffer;
  uartCtrl_1 : entity work.UartCtrl
    port map ( 
      io_config_frame_dataLength => bridge_uartConfigReg_frame_dataLength,
      io_config_frame_stop => bridge_uartConfigReg_frame_stop,
      io_config_frame_parity => bridge_uartConfigReg_frame_parity,
      io_config_clockDivider => bridge_uartConfigReg_clockDivider,
      io_write_valid => bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid,
      io_write_ready => uartCtrl_1_io_write_ready,
      io_write_payload => bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_payload,
      io_read_valid => uartCtrl_1_io_read_valid,
      io_read_ready => uartCtrl_1_io_read_queueWithOccupancy_io_push_ready,
      io_read_payload => uartCtrl_1_io_read_payload,
      io_uart_txd => uartCtrl_1_io_uart_txd,
      io_uart_rxd => io_uart_rxd,
      io_readError => uartCtrl_1_io_readError,
      io_writeBreak => bridge_misc_doBreak,
      io_readBreak => uartCtrl_1_io_readBreak,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  bridge_write_streamUnbuffered_queueWithOccupancy : entity work.StreamFifo
    port map ( 
      io_push_valid => bridge_write_streamUnbuffered_valid,
      io_push_ready => bridge_write_streamUnbuffered_queueWithOccupancy_io_push_ready,
      io_push_payload => bridge_write_streamUnbuffered_payload,
      io_pop_valid => bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid,
      io_pop_ready => uartCtrl_1_io_write_ready,
      io_pop_payload => bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_payload,
      io_flush => pkg_toStdLogic(false),
      io_occupancy => bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy,
      io_availability => bridge_write_streamUnbuffered_queueWithOccupancy_io_availability,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  uartCtrl_1_io_read_queueWithOccupancy : entity work.StreamFifo
    port map ( 
      io_push_valid => uartCtrl_1_io_read_valid,
      io_push_ready => uartCtrl_1_io_read_queueWithOccupancy_io_push_ready,
      io_push_payload => uartCtrl_1_io_read_payload,
      io_pop_valid => uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid,
      io_pop_ready => uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready,
      io_pop_payload => uartCtrl_1_io_read_queueWithOccupancy_io_pop_payload,
      io_flush => pkg_toStdLogic(false),
      io_occupancy => uartCtrl_1_io_read_queueWithOccupancy_io_occupancy,
      io_availability => uartCtrl_1_io_read_queueWithOccupancy_io_availability,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  io_uart_txd <= uartCtrl_1_io_uart_txd;
  io_apb_PREADY_read_buffer <= pkg_toStdLogic(true);
  process(io_apb_PADDR,bridge_read_streamBreaked_valid,bridge_read_streamBreaked_payload,bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy,bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid,uartCtrl_1_io_read_queueWithOccupancy_io_occupancy,bridge_interruptCtrl_writeIntEnable,bridge_interruptCtrl_readIntEnable,bridge_interruptCtrl_writeInt,bridge_interruptCtrl_readInt,bridge_misc_readError,bridge_misc_readOverflowError,uartCtrl_1_io_readBreak,bridge_misc_breakDetected)
  begin
    io_apb_PRDATA <= pkg_stdLogicVector("00000000000000000000000000000000");
    case io_apb_PADDR is
      when "00000" =>
        io_apb_PRDATA(16 downto 16) <= pkg_toStdLogicVector((bridge_read_streamBreaked_valid xor pkg_toStdLogic(false)));
        io_apb_PRDATA(7 downto 0) <= bridge_read_streamBreaked_payload;
      when "00100" =>
        io_apb_PRDATA(20 downto 16) <= std_logic_vector((pkg_unsigned("10000") - bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy));
        io_apb_PRDATA(15 downto 15) <= pkg_toStdLogicVector(bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid);
        io_apb_PRDATA(28 downto 24) <= std_logic_vector(uartCtrl_1_io_read_queueWithOccupancy_io_occupancy);
        io_apb_PRDATA(0 downto 0) <= pkg_toStdLogicVector(bridge_interruptCtrl_writeIntEnable);
        io_apb_PRDATA(1 downto 1) <= pkg_toStdLogicVector(bridge_interruptCtrl_readIntEnable);
        io_apb_PRDATA(8 downto 8) <= pkg_toStdLogicVector(bridge_interruptCtrl_writeInt);
        io_apb_PRDATA(9 downto 9) <= pkg_toStdLogicVector(bridge_interruptCtrl_readInt);
      when "10000" =>
        io_apb_PRDATA(0 downto 0) <= pkg_toStdLogicVector(bridge_misc_readError);
        io_apb_PRDATA(1 downto 1) <= pkg_toStdLogicVector(bridge_misc_readOverflowError);
        io_apb_PRDATA(8 downto 8) <= pkg_toStdLogicVector(uartCtrl_1_io_readBreak);
        io_apb_PRDATA(9 downto 9) <= pkg_toStdLogicVector(bridge_misc_breakDetected);
      when others =>
    end case;
  end process;

  busCtrl_askWrite <= ((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PWRITE);
  busCtrl_askRead <= ((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and (not io_apb_PWRITE));
  busCtrl_doWrite <= (((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PREADY_read_buffer) and io_apb_PWRITE);
  busCtrl_doRead <= (((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PREADY_read_buffer) and (not io_apb_PWRITE));
  bridge_uartConfigReg_clockDivider <= zz_bridge_uartConfigReg_clockDivider;
  bridge_uartConfigReg_frame_dataLength <= pkg_unsigned("111");
  bridge_uartConfigReg_frame_parity <= UartParityType_seq_NONE;
  bridge_uartConfigReg_frame_stop <= UartStopType_seq_ONE;
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    zz_bridge_write_streamUnbuffered_valid <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "00000" =>
        if busCtrl_doWrite = '1' then
          zz_bridge_write_streamUnbuffered_valid <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  bridge_write_streamUnbuffered_valid <= zz_bridge_write_streamUnbuffered_valid;
  bridge_write_streamUnbuffered_payload <= pkg_extract(io_apb_PWDATA,7,0);
  bridge_write_streamUnbuffered_ready <= bridge_write_streamUnbuffered_queueWithOccupancy_io_push_ready;
  process(uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid,uartCtrl_1_io_readBreak)
  begin
    bridge_read_streamBreaked_valid <= uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid;
    if uartCtrl_1_io_readBreak = '1' then
      bridge_read_streamBreaked_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  process(bridge_read_streamBreaked_ready,uartCtrl_1_io_readBreak)
  begin
    uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready <= bridge_read_streamBreaked_ready;
    if uartCtrl_1_io_readBreak = '1' then
      uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  bridge_read_streamBreaked_payload <= uartCtrl_1_io_read_queueWithOccupancy_io_pop_payload;
  process(io_apb_PADDR,busCtrl_doRead)
  begin
    bridge_read_streamBreaked_ready <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "00000" =>
        if busCtrl_doRead = '1' then
          bridge_read_streamBreaked_ready <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  bridge_interruptCtrl_readInt <= (bridge_interruptCtrl_readIntEnable and bridge_read_streamBreaked_valid);
  bridge_interruptCtrl_writeInt <= (bridge_interruptCtrl_writeIntEnable and (not bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid));
  bridge_interruptCtrl_interrupt <= (bridge_interruptCtrl_readInt or bridge_interruptCtrl_writeInt);
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_BusSlaveFactory_l335 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "10000" =>
        if busCtrl_doWrite = '1' then
          when_BusSlaveFactory_l335 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  when_BusSlaveFactory_l337 <= pkg_extract(io_apb_PWDATA,0);
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_BusSlaveFactory_l335_1 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "10000" =>
        if busCtrl_doWrite = '1' then
          when_BusSlaveFactory_l335_1 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  when_BusSlaveFactory_l337_1 <= pkg_extract(io_apb_PWDATA,1);
  uartCtrl_1_io_read_isStall <= (uartCtrl_1_io_read_valid and (not uartCtrl_1_io_read_queueWithOccupancy_io_push_ready));
  when_UartCtrl_l155 <= (uartCtrl_1_io_readBreak and (not uartCtrl_1_io_readBreak_regNext));
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_BusSlaveFactory_l335_2 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "10000" =>
        if busCtrl_doWrite = '1' then
          when_BusSlaveFactory_l335_2 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  when_BusSlaveFactory_l337_2 <= pkg_extract(io_apb_PWDATA,9);
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_BusSlaveFactory_l366 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "10000" =>
        if busCtrl_doWrite = '1' then
          when_BusSlaveFactory_l366 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  when_BusSlaveFactory_l368 <= pkg_extract(io_apb_PWDATA,10);
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_BusSlaveFactory_l335_3 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "10000" =>
        if busCtrl_doWrite = '1' then
          when_BusSlaveFactory_l335_3 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  when_BusSlaveFactory_l337_3 <= pkg_extract(io_apb_PWDATA,11);
  io_interrupt <= bridge_interruptCtrl_interrupt;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      bridge_interruptCtrl_writeIntEnable <= pkg_toStdLogic(false);
      bridge_interruptCtrl_readIntEnable <= pkg_toStdLogic(false);
      bridge_misc_readError <= pkg_toStdLogic(false);
      bridge_misc_readOverflowError <= pkg_toStdLogic(false);
      bridge_misc_breakDetected <= pkg_toStdLogic(false);
      bridge_misc_doBreak <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if when_BusSlaveFactory_l335 = '1' then
        if when_BusSlaveFactory_l337 = '1' then
          bridge_misc_readError <= pkg_extract(pkg_stdLogicVector("0"),0);
        end if;
      end if;
      if uartCtrl_1_io_readError = '1' then
        bridge_misc_readError <= pkg_toStdLogic(true);
      end if;
      if when_BusSlaveFactory_l335_1 = '1' then
        if when_BusSlaveFactory_l337_1 = '1' then
          bridge_misc_readOverflowError <= pkg_extract(pkg_stdLogicVector("0"),0);
        end if;
      end if;
      if uartCtrl_1_io_read_isStall = '1' then
        bridge_misc_readOverflowError <= pkg_toStdLogic(true);
      end if;
      if when_UartCtrl_l155 = '1' then
        bridge_misc_breakDetected <= pkg_toStdLogic(true);
      end if;
      if when_BusSlaveFactory_l335_2 = '1' then
        if when_BusSlaveFactory_l337_2 = '1' then
          bridge_misc_breakDetected <= pkg_extract(pkg_stdLogicVector("0"),0);
        end if;
      end if;
      if when_BusSlaveFactory_l366 = '1' then
        if when_BusSlaveFactory_l368 = '1' then
          bridge_misc_doBreak <= pkg_extract(pkg_stdLogicVector("1"),0);
        end if;
      end if;
      if when_BusSlaveFactory_l335_3 = '1' then
        if when_BusSlaveFactory_l337_3 = '1' then
          bridge_misc_doBreak <= pkg_extract(pkg_stdLogicVector("0"),0);
        end if;
      end if;
      case io_apb_PADDR is
        when "00100" =>
          if busCtrl_doWrite = '1' then
            bridge_interruptCtrl_writeIntEnable <= pkg_extract(io_apb_PWDATA,0);
            bridge_interruptCtrl_readIntEnable <= pkg_extract(io_apb_PWDATA,1);
          end if;
        when others =>
      end case;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      uartCtrl_1_io_readBreak_regNext <= uartCtrl_1_io_readBreak;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity MuraxApb3Timer is
  port(
    io_apb_PADDR : in unsigned(7 downto 0);
    io_apb_PSEL : in std_logic_vector(0 downto 0);
    io_apb_PENABLE : in std_logic;
    io_apb_PREADY : out std_logic;
    io_apb_PWRITE : in std_logic;
    io_apb_PWDATA : in std_logic_vector(31 downto 0);
    io_apb_PRDATA : out std_logic_vector(31 downto 0);
    io_apb_PSLVERROR : out std_logic;
    io_interrupt : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end MuraxApb3Timer;

architecture arch of MuraxApb3Timer is
  signal timerA_io_tick : std_logic;
  signal timerA_io_clear : std_logic;
  signal timerB_io_tick : std_logic;
  signal timerB_io_clear : std_logic;
  signal interruptCtrl_1_io_inputs : std_logic_vector(1 downto 0);
  signal interruptCtrl_1_io_clears : std_logic_vector(1 downto 0);
  signal io_apb_PREADY_read_buffer : std_logic;
  signal prescaler_1_io_overflow : std_logic;
  signal timerA_io_full : std_logic;
  signal timerA_io_value : unsigned(15 downto 0);
  signal timerB_io_full : std_logic;
  signal timerB_io_value : unsigned(15 downto 0);
  signal interruptCtrl_1_io_pendings : std_logic_vector(1 downto 0);

  signal busCtrl_askWrite : std_logic;
  signal busCtrl_askRead : std_logic;
  signal busCtrl_doWrite : std_logic;
  signal busCtrl_doRead : std_logic;
  signal zz_io_limit : unsigned(31 downto 0);
  signal zz_io_clear : std_logic;
  signal timerABridge_ticksEnable : std_logic_vector(1 downto 0);
  signal timerABridge_clearsEnable : std_logic_vector(0 downto 0);
  signal timerABridge_busClearing : std_logic;
  signal timerA_io_limit_driver : unsigned(15 downto 0);
  signal when_Timer_l40 : std_logic;
  signal when_Timer_l44 : std_logic;
  signal timerBBridge_ticksEnable : std_logic_vector(1 downto 0);
  signal timerBBridge_clearsEnable : std_logic_vector(0 downto 0);
  signal timerBBridge_busClearing : std_logic;
  signal timerB_io_limit_driver : unsigned(15 downto 0);
  signal when_Timer_l40_1 : std_logic;
  signal when_Timer_l44_1 : std_logic;
  signal interruptCtrl_1_io_masks_driver : std_logic_vector(1 downto 0);
begin
  io_apb_PREADY <= io_apb_PREADY_read_buffer;
  prescaler_1 : entity work.Prescaler
    port map ( 
      io_clear => zz_io_clear,
      io_limit => zz_io_limit,
      io_overflow => prescaler_1_io_overflow,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  timerA : entity work.Timer
    port map ( 
      io_tick => timerA_io_tick,
      io_clear => timerA_io_clear,
      io_limit => timerA_io_limit_driver,
      io_full => timerA_io_full,
      io_value => timerA_io_value,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  timerB : entity work.Timer
    port map ( 
      io_tick => timerB_io_tick,
      io_clear => timerB_io_clear,
      io_limit => timerB_io_limit_driver,
      io_full => timerB_io_full,
      io_value => timerB_io_value,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  interruptCtrl_1 : entity work.InterruptCtrl
    port map ( 
      io_inputs => interruptCtrl_1_io_inputs,
      io_clears => interruptCtrl_1_io_clears,
      io_masks => interruptCtrl_1_io_masks_driver,
      io_pendings => interruptCtrl_1_io_pendings,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  io_apb_PREADY_read_buffer <= pkg_toStdLogic(true);
  process(io_apb_PADDR,zz_io_limit,timerABridge_ticksEnable,timerABridge_clearsEnable,timerA_io_limit_driver,timerA_io_value,timerBBridge_ticksEnable,timerBBridge_clearsEnable,timerB_io_limit_driver,timerB_io_value,interruptCtrl_1_io_pendings,interruptCtrl_1_io_masks_driver)
  begin
    io_apb_PRDATA <= pkg_stdLogicVector("00000000000000000000000000000000");
    case io_apb_PADDR is
      when "00000000" =>
        io_apb_PRDATA(31 downto 0) <= std_logic_vector(zz_io_limit);
      when "01000000" =>
        io_apb_PRDATA(1 downto 0) <= timerABridge_ticksEnable;
        io_apb_PRDATA(16 downto 16) <= timerABridge_clearsEnable;
      when "01000100" =>
        io_apb_PRDATA(15 downto 0) <= std_logic_vector(timerA_io_limit_driver);
      when "01001000" =>
        io_apb_PRDATA(15 downto 0) <= std_logic_vector(timerA_io_value);
      when "01010000" =>
        io_apb_PRDATA(1 downto 0) <= timerBBridge_ticksEnable;
        io_apb_PRDATA(16 downto 16) <= timerBBridge_clearsEnable;
      when "01010100" =>
        io_apb_PRDATA(15 downto 0) <= std_logic_vector(timerB_io_limit_driver);
      when "01011000" =>
        io_apb_PRDATA(15 downto 0) <= std_logic_vector(timerB_io_value);
      when "00010000" =>
        io_apb_PRDATA(1 downto 0) <= interruptCtrl_1_io_pendings;
      when "00010100" =>
        io_apb_PRDATA(1 downto 0) <= interruptCtrl_1_io_masks_driver;
      when others =>
    end case;
  end process;

  io_apb_PSLVERROR <= pkg_toStdLogic(false);
  busCtrl_askWrite <= ((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PWRITE);
  busCtrl_askRead <= ((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and (not io_apb_PWRITE));
  busCtrl_doWrite <= (((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PREADY_read_buffer) and io_apb_PWRITE);
  busCtrl_doRead <= (((pkg_extract(io_apb_PSEL,0) and io_apb_PENABLE) and io_apb_PREADY_read_buffer) and (not io_apb_PWRITE));
  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    zz_io_clear <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "00000000" =>
        if busCtrl_doWrite = '1' then
          zz_io_clear <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  process(when_Timer_l40,when_Timer_l44)
  begin
    timerABridge_busClearing <= pkg_toStdLogic(false);
    if when_Timer_l40 = '1' then
      timerABridge_busClearing <= pkg_toStdLogic(true);
    end if;
    if when_Timer_l44 = '1' then
      timerABridge_busClearing <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_Timer_l40 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "01000100" =>
        if busCtrl_doWrite = '1' then
          when_Timer_l40 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_Timer_l44 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "01001000" =>
        if busCtrl_doWrite = '1' then
          when_Timer_l44 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  timerA_io_clear <= (pkg_toStdLogic((timerABridge_clearsEnable and pkg_toStdLogicVector(timerA_io_full)) /= pkg_stdLogicVector("0")) or timerABridge_busClearing);
  timerA_io_tick <= pkg_toStdLogic((timerABridge_ticksEnable and pkg_cat(pkg_toStdLogicVector(prescaler_1_io_overflow),pkg_toStdLogicVector(pkg_toStdLogic(true)))) /= pkg_stdLogicVector("00"));
  process(when_Timer_l40_1,when_Timer_l44_1)
  begin
    timerBBridge_busClearing <= pkg_toStdLogic(false);
    if when_Timer_l40_1 = '1' then
      timerBBridge_busClearing <= pkg_toStdLogic(true);
    end if;
    if when_Timer_l44_1 = '1' then
      timerBBridge_busClearing <= pkg_toStdLogic(true);
    end if;
  end process;

  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_Timer_l40_1 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "01010100" =>
        if busCtrl_doWrite = '1' then
          when_Timer_l40_1 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  process(io_apb_PADDR,busCtrl_doWrite)
  begin
    when_Timer_l44_1 <= pkg_toStdLogic(false);
    case io_apb_PADDR is
      when "01011000" =>
        if busCtrl_doWrite = '1' then
          when_Timer_l44_1 <= pkg_toStdLogic(true);
        end if;
      when others =>
    end case;
  end process;

  timerB_io_clear <= (pkg_toStdLogic((timerBBridge_clearsEnable and pkg_toStdLogicVector(timerB_io_full)) /= pkg_stdLogicVector("0")) or timerBBridge_busClearing);
  timerB_io_tick <= pkg_toStdLogic((timerBBridge_ticksEnable and pkg_cat(pkg_toStdLogicVector(prescaler_1_io_overflow),pkg_toStdLogicVector(pkg_toStdLogic(true)))) /= pkg_stdLogicVector("00"));
  process(io_apb_PADDR,busCtrl_doWrite,io_apb_PWDATA)
  begin
    interruptCtrl_1_io_clears <= pkg_stdLogicVector("00");
    case io_apb_PADDR is
      when "00010000" =>
        if busCtrl_doWrite = '1' then
          interruptCtrl_1_io_clears <= pkg_extract(io_apb_PWDATA,1,0);
        end if;
      when others =>
    end case;
  end process;

  process(timerA_io_full,timerB_io_full)
  begin
    interruptCtrl_1_io_inputs(0) <= timerA_io_full;
    interruptCtrl_1_io_inputs(1) <= timerB_io_full;
  end process;

  io_interrupt <= pkg_toStdLogic(interruptCtrl_1_io_pendings /= pkg_stdLogicVector("00"));
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      timerABridge_ticksEnable <= pkg_stdLogicVector("00");
      timerABridge_clearsEnable <= pkg_stdLogicVector("0");
      timerBBridge_ticksEnable <= pkg_stdLogicVector("00");
      timerBBridge_clearsEnable <= pkg_stdLogicVector("0");
      interruptCtrl_1_io_masks_driver <= pkg_stdLogicVector("00");
    elsif rising_edge(io_mainClk) then
      case io_apb_PADDR is
        when "01000000" =>
          if busCtrl_doWrite = '1' then
            timerABridge_ticksEnable <= pkg_extract(io_apb_PWDATA,1,0);
            timerABridge_clearsEnable <= pkg_extract(io_apb_PWDATA,16,16);
          end if;
        when "01010000" =>
          if busCtrl_doWrite = '1' then
            timerBBridge_ticksEnable <= pkg_extract(io_apb_PWDATA,1,0);
            timerBBridge_clearsEnable <= pkg_extract(io_apb_PWDATA,16,16);
          end if;
        when "00010100" =>
          if busCtrl_doWrite = '1' then
            interruptCtrl_1_io_masks_driver <= pkg_extract(io_apb_PWDATA,1,0);
          end if;
        when others =>
      end case;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      case io_apb_PADDR is
        when "00000000" =>
          if busCtrl_doWrite = '1' then
            zz_io_limit <= unsigned(pkg_extract(io_apb_PWDATA,31,0));
          end if;
        when "01000100" =>
          if busCtrl_doWrite = '1' then
            timerA_io_limit_driver <= unsigned(pkg_extract(io_apb_PWDATA,15,0));
          end if;
        when "01010100" =>
          if busCtrl_doWrite = '1' then
            timerB_io_limit_driver <= unsigned(pkg_extract(io_apb_PWDATA,15,0));
          end if;
        when others =>
      end case;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity VexRiscv is
  port(
    dBus_cmd_valid : out std_logic;
    dBus_cmd_ready : in std_logic;
    dBus_cmd_payload_wr : out std_logic;
    dBus_cmd_payload_uncached : out std_logic;
    dBus_cmd_payload_address : out unsigned(31 downto 0);
    dBus_cmd_payload_data : out std_logic_vector(31 downto 0);
    dBus_cmd_payload_mask : out std_logic_vector(3 downto 0);
    dBus_cmd_payload_size : out unsigned(2 downto 0);
    dBus_cmd_payload_last : out std_logic;
    dBus_rsp_valid : in std_logic;
    dBus_rsp_payload_last : in std_logic;
    dBus_rsp_payload_data : in std_logic_vector(31 downto 0);
    dBus_rsp_payload_error : in std_logic;
    timerInterrupt : in std_logic;
    externalInterrupt : in std_logic;
    softwareInterrupt : in std_logic;
    debug_bus_cmd_valid : in std_logic;
    debug_bus_cmd_ready : out std_logic;
    debug_bus_cmd_payload_wr : in std_logic;
    debug_bus_cmd_payload_address : in unsigned(7 downto 0);
    debug_bus_cmd_payload_data : in std_logic_vector(31 downto 0);
    debug_bus_rsp_data : out std_logic_vector(31 downto 0);
    debug_resetOut : out std_logic;
    iBus_cmd_valid : out std_logic;
    iBus_cmd_ready : in std_logic;
    iBus_cmd_payload_address : out unsigned(31 downto 0);
    iBus_cmd_payload_size : out unsigned(2 downto 0);
    iBus_rsp_valid : in std_logic;
    iBus_rsp_payload_data : in std_logic_vector(31 downto 0);
    iBus_rsp_payload_error : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic;
    resetCtrl_systemReset : in std_logic
  );
end VexRiscv;

architecture arch of VexRiscv is
  signal IBusCachedPlugin_cache_io_flush : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_prefetch_isValid : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_fetch_isValid : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_fetch_isStuck : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_fetch_isRemoved : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_isValid : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_isStuck : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_isUser : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_fill_valid : std_logic;
  signal dataCache_1_io_cpu_execute_isValid : std_logic;
  signal dataCache_1_io_cpu_execute_address : unsigned(31 downto 0);
  signal dataCache_1_io_cpu_memory_isValid : std_logic;
  signal dataCache_1_io_cpu_memory_address : unsigned(31 downto 0);
  signal dataCache_1_io_cpu_memory_mmuRsp_isIoAccess : std_logic;
  signal dataCache_1_io_cpu_writeBack_isValid : std_logic;
  signal dataCache_1_io_cpu_writeBack_isUser : std_logic;
  signal dataCache_1_io_cpu_writeBack_storeData : std_logic_vector(31 downto 0);
  signal dataCache_1_io_cpu_writeBack_address : unsigned(31 downto 0);
  signal dataCache_1_io_cpu_writeBack_fence_SW : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_SR : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_SO : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_SI : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_PW : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_PR : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_PO : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_PI : std_logic;
  signal dataCache_1_io_cpu_writeBack_fence_FM : std_logic_vector(3 downto 0);
  signal dataCache_1_io_cpu_flush_valid : std_logic;
  signal zz_IBusCachedPlugin_predictor_history_port0 : std_logic_vector(55 downto 0);
  signal zz_RegFilePlugin_regFile_port0 : std_logic_vector(31 downto 0);
  signal zz_RegFilePlugin_regFile_port0_1 : std_logic_vector(31 downto 0);
  signal debug_bus_cmd_ready_read_buffer : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_prefetch_haltIt : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_fetch_data : std_logic_vector(31 downto 0);
  signal IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress : unsigned(31 downto 0);
  signal IBusCachedPlugin_cache_io_cpu_decode_error : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_mmuException : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_data : std_logic_vector(31 downto 0);
  signal IBusCachedPlugin_cache_io_cpu_decode_cacheMiss : std_logic;
  signal IBusCachedPlugin_cache_io_cpu_decode_physicalAddress : unsigned(31 downto 0);
  signal IBusCachedPlugin_cache_io_mem_cmd_valid : std_logic;
  signal IBusCachedPlugin_cache_io_mem_cmd_payload_address : unsigned(31 downto 0);
  signal IBusCachedPlugin_cache_io_mem_cmd_payload_size : unsigned(2 downto 0);
  signal dataCache_1_io_cpu_execute_haltIt : std_logic;
  signal dataCache_1_io_cpu_execute_refilling : std_logic;
  signal dataCache_1_io_cpu_memory_isWrite : std_logic;
  signal dataCache_1_io_cpu_writeBack_haltIt : std_logic;
  signal dataCache_1_io_cpu_writeBack_data : std_logic_vector(31 downto 0);
  signal dataCache_1_io_cpu_writeBack_mmuException : std_logic;
  signal dataCache_1_io_cpu_writeBack_unalignedAccess : std_logic;
  signal dataCache_1_io_cpu_writeBack_accessError : std_logic;
  signal dataCache_1_io_cpu_writeBack_isWrite : std_logic;
  signal dataCache_1_io_cpu_writeBack_keepMemRspData : std_logic;
  signal dataCache_1_io_cpu_writeBack_exclusiveOk : std_logic;
  signal dataCache_1_io_cpu_flush_ready : std_logic;
  signal dataCache_1_io_cpu_redo : std_logic;
  signal dataCache_1_io_mem_cmd_valid : std_logic;
  signal dataCache_1_io_mem_cmd_payload_wr : std_logic;
  signal dataCache_1_io_mem_cmd_payload_uncached : std_logic;
  signal dataCache_1_io_mem_cmd_payload_address : unsigned(31 downto 0);
  signal dataCache_1_io_mem_cmd_payload_data : std_logic_vector(31 downto 0);
  signal dataCache_1_io_mem_cmd_payload_mask : std_logic_vector(3 downto 0);
  signal dataCache_1_io_mem_cmd_payload_size : unsigned(2 downto 0);
  signal dataCache_1_io_mem_cmd_payload_last : std_logic;
  signal zz_decode_LEGAL_INSTRUCTION : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_1 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_2 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_3 : std_logic;
  signal zz_decode_LEGAL_INSTRUCTION_4 : std_logic_vector(0 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_5 : std_logic_vector(13 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_6 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_7 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_8 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_9 : std_logic;
  signal zz_decode_LEGAL_INSTRUCTION_10 : std_logic_vector(0 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_11 : std_logic_vector(7 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_12 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_13 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_14 : std_logic_vector(31 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_15 : std_logic;
  signal zz_decode_LEGAL_INSTRUCTION_16 : std_logic_vector(0 downto 0);
  signal zz_decode_LEGAL_INSTRUCTION_17 : std_logic_vector(1 downto 0);
  signal zz_IBusCachedPlugin_jump_pcLoad_payload_4 : unsigned(31 downto 0);
  signal zz_IBusCachedPlugin_jump_pcLoad_payload_5 : unsigned(1 downto 0);
  signal zz_IBusCachedPlugin_predictor_history_port : std_logic_vector(55 downto 0);
  signal zz_IBusCachedPlugin_predictor_history_port_1 : unsigned(7 downto 0);
  signal zz_zz_IBusCachedPlugin_predictor_buffer_line_source_1 : unsigned(7 downto 0);
  signal zz_writeBack_DBusCachedPlugin_rspShifted : std_logic_vector(7 downto 0);
  signal zz_writeBack_DBusCachedPlugin_rspShifted_1 : unsigned(1 downto 0);
  signal zz_writeBack_DBusCachedPlugin_rspShifted_2 : std_logic_vector(7 downto 0);
  signal zz_writeBack_DBusCachedPlugin_rspShifted_3 : unsigned(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_1 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_2 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_3 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_4 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_5 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_6 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_7 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_8 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_9 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_10 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_11 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_12 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_13 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_14 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_15 : std_logic_vector(25 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_16 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_17 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_18 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_19 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_20 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_21 : std_logic_vector(22 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_22 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_23 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_24 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_25 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_26 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_27 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_28 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_29 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_30 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_31 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_32 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_33 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_34 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_35 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_36 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_37 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_38 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_39 : std_logic_vector(17 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_40 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_41 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_42 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_43 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_44 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_45 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_46 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_47 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_48 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_49 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_50 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_51 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_52 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_53 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_54 : std_logic_vector(14 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_55 : std_logic_vector(2 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_56 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_57 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_58 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_59 : std_logic_vector(2 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_60 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_61 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_62 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_63 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_64 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_65 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_66 : std_logic_vector(3 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_67 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_68 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_69 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_70 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_71 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_72 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_73 : std_logic_vector(11 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_74 : std_logic_vector(2 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_75 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_76 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_77 : std_logic_vector(2 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_78 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_79 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_80 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_81 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_82 : std_logic_vector(3 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_83 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_84 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_85 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_86 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_87 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_88 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_89 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_90 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_91 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_92 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_93 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_94 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_95 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_96 : std_logic_vector(8 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_97 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_98 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_99 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_100 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_101 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_102 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_103 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_104 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_105 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_106 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_107 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_108 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_109 : std_logic_vector(5 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_110 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_111 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_112 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_113 : std_logic_vector(2 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_114 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_115 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_116 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_117 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_118 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_119 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_120 : std_logic_vector(3 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_121 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_122 : std_logic;
  signal zz_zz_decode_ENV_CTRL_2_123 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_124 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_125 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_126 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_127 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_128 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_129 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_130 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_131 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_132 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_133 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_134 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_135 : std_logic_vector(1 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_136 : std_logic_vector(0 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_137 : std_logic_vector(31 downto 0);
  signal zz_zz_decode_ENV_CTRL_2_138 : std_logic_vector(0 downto 0);
  signal zz_RegFilePlugin_regFile_port : std_logic;
  signal zz_decode_RegFilePlugin_rs1Data : std_logic;
  signal zz_RegFilePlugin_regFile_port_1 : std_logic;
  signal zz_decode_RegFilePlugin_rs2Data : std_logic;
  signal zz_when : std_logic;
  attribute keep : boolean;
  attribute syn_keep : boolean;

  signal memory_MUL_LOW : signed(51 downto 0);
  signal execute_TARGET_MISSMATCH2 : std_logic;
  signal execute_NEXT_PC2 : unsigned(31 downto 0);
  signal execute_BRANCH_DO : std_logic;
  signal memory_MUL_HH : signed(33 downto 0);
  signal execute_MUL_HH : signed(33 downto 0);
  signal execute_MUL_HL : signed(33 downto 0);
  signal execute_MUL_LH : signed(33 downto 0);
  signal execute_MUL_LL : unsigned(31 downto 0);
  signal execute_REGFILE_WRITE_DATA : std_logic_vector(31 downto 0);
  signal memory_MEMORY_STORE_DATA_RF : std_logic_vector(31 downto 0);
  signal execute_MEMORY_STORE_DATA_RF : std_logic_vector(31 downto 0);
  signal decode_DO_EBREAK : std_logic;
  signal decode_CSR_READ_OPCODE : std_logic;
  signal decode_CSR_WRITE_OPCODE : std_logic;
  signal decode_SRC2_FORCE_ZERO : std_logic;
  signal zz_memory_to_writeBack_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_memory_to_writeBack_ENV_CTRL_1 : EnvCtrlEnum_seq_type;
  signal zz_execute_to_memory_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_execute_to_memory_ENV_CTRL_1 : EnvCtrlEnum_seq_type;
  signal decode_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_decode_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_decode_to_execute_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_decode_to_execute_ENV_CTRL_1 : EnvCtrlEnum_seq_type;
  signal decode_IS_CSR : std_logic;
  signal decode_BRANCH_CTRL : BranchCtrlEnum_seq_type;
  signal zz_decode_BRANCH_CTRL : BranchCtrlEnum_seq_type;
  signal zz_decode_to_execute_BRANCH_CTRL : BranchCtrlEnum_seq_type;
  signal zz_decode_to_execute_BRANCH_CTRL_1 : BranchCtrlEnum_seq_type;
  signal decode_IS_RS2_SIGNED : std_logic;
  signal decode_IS_RS1_SIGNED : std_logic;
  signal decode_IS_DIV : std_logic;
  signal memory_IS_MUL : std_logic;
  signal execute_IS_MUL : std_logic;
  signal decode_IS_MUL : std_logic;
  signal decode_SHIFT_CTRL : ShiftCtrlEnum_seq_type;
  signal zz_decode_SHIFT_CTRL : ShiftCtrlEnum_seq_type;
  signal zz_decode_to_execute_SHIFT_CTRL : ShiftCtrlEnum_seq_type;
  signal zz_decode_to_execute_SHIFT_CTRL_1 : ShiftCtrlEnum_seq_type;
  signal decode_ALU_BITWISE_CTRL : AluBitwiseCtrlEnum_seq_type;
  signal zz_decode_ALU_BITWISE_CTRL : AluBitwiseCtrlEnum_seq_type;
  signal zz_decode_to_execute_ALU_BITWISE_CTRL : AluBitwiseCtrlEnum_seq_type;
  signal zz_decode_to_execute_ALU_BITWISE_CTRL_1 : AluBitwiseCtrlEnum_seq_type;
  signal decode_SRC_LESS_UNSIGNED : std_logic;
  signal decode_MEMORY_MANAGMENT : std_logic;
  signal memory_MEMORY_WR : std_logic;
  signal decode_MEMORY_WR : std_logic;
  signal execute_BYPASSABLE_MEMORY_STAGE : std_logic;
  signal decode_BYPASSABLE_MEMORY_STAGE : std_logic;
  signal decode_BYPASSABLE_EXECUTE_STAGE : std_logic;
  signal decode_SRC2_CTRL : Src2CtrlEnum_seq_type;
  signal zz_decode_SRC2_CTRL : Src2CtrlEnum_seq_type;
  signal zz_decode_to_execute_SRC2_CTRL : Src2CtrlEnum_seq_type;
  signal zz_decode_to_execute_SRC2_CTRL_1 : Src2CtrlEnum_seq_type;
  signal decode_ALU_CTRL : AluCtrlEnum_seq_type;
  signal zz_decode_ALU_CTRL : AluCtrlEnum_seq_type;
  signal zz_decode_to_execute_ALU_CTRL : AluCtrlEnum_seq_type;
  signal zz_decode_to_execute_ALU_CTRL_1 : AluCtrlEnum_seq_type;
  signal decode_SRC1_CTRL : Src1CtrlEnum_seq_type;
  signal zz_decode_SRC1_CTRL : Src1CtrlEnum_seq_type;
  signal zz_decode_to_execute_SRC1_CTRL : Src1CtrlEnum_seq_type;
  signal zz_decode_to_execute_SRC1_CTRL_1 : Src1CtrlEnum_seq_type;
  signal decode_MEMORY_FORCE_CONSTISTENCY : std_logic;
  signal execute_PREDICTION_CONTEXT_hazard : std_logic;
  signal execute_PREDICTION_CONTEXT_hit : std_logic;
  signal execute_PREDICTION_CONTEXT_line_source : std_logic_vector(21 downto 0);
  signal execute_PREDICTION_CONTEXT_line_branchWish : unsigned(1 downto 0);
  signal execute_PREDICTION_CONTEXT_line_target : unsigned(31 downto 0);
  signal decode_PREDICTION_CONTEXT_hazard : std_logic;
  signal decode_PREDICTION_CONTEXT_hit : std_logic;
  signal decode_PREDICTION_CONTEXT_line_source : std_logic_vector(21 downto 0);
  signal decode_PREDICTION_CONTEXT_line_branchWish : unsigned(1 downto 0);
  signal decode_PREDICTION_CONTEXT_line_target : unsigned(31 downto 0);
  signal writeBack_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal memory_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal execute_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal decode_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal execute_DO_EBREAK : std_logic;
  signal decode_IS_EBREAK : std_logic;
  signal execute_CSR_READ_OPCODE : std_logic;
  signal execute_CSR_WRITE_OPCODE : std_logic;
  signal execute_IS_CSR : std_logic;
  signal memory_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_memory_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal execute_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_execute_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal writeBack_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal zz_writeBack_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal memory_NEXT_PC2 : unsigned(31 downto 0);
  signal memory_PC : unsigned(31 downto 0);
  signal memory_BRANCH_CALC : unsigned(31 downto 0);
  signal memory_TARGET_MISSMATCH2 : std_logic;
  signal memory_BRANCH_DO : std_logic;
  signal execute_BRANCH_CALC : unsigned(31 downto 0);
  signal execute_BRANCH_SRC22 : unsigned(31 downto 0);
  signal execute_PC : unsigned(31 downto 0);
  signal execute_BRANCH_CTRL : BranchCtrlEnum_seq_type;
  signal zz_execute_BRANCH_CTRL : BranchCtrlEnum_seq_type;
  signal decode_RS2_USE : std_logic;
  signal decode_RS1_USE : std_logic;
  signal execute_REGFILE_WRITE_VALID : std_logic;
  signal execute_BYPASSABLE_EXECUTE_STAGE : std_logic;
  signal memory_REGFILE_WRITE_VALID : std_logic;
  signal memory_BYPASSABLE_MEMORY_STAGE : std_logic;
  signal writeBack_REGFILE_WRITE_VALID : std_logic;
  signal decode_RS2 : std_logic_vector(31 downto 0);
  signal decode_RS1 : std_logic_vector(31 downto 0);
  signal execute_IS_RS1_SIGNED : std_logic;
  signal execute_IS_DIV : std_logic;
  signal execute_IS_RS2_SIGNED : std_logic;
  signal zz_decode_RS2 : std_logic_vector(31 downto 0);
  signal memory_INSTRUCTION : std_logic_vector(31 downto 0);
  signal memory_IS_DIV : std_logic;
  signal writeBack_IS_MUL : std_logic;
  signal writeBack_MUL_HH : signed(33 downto 0);
  signal writeBack_MUL_LOW : signed(51 downto 0);
  signal memory_MUL_HL : signed(33 downto 0);
  signal memory_MUL_LH : signed(33 downto 0);
  signal memory_MUL_LL : unsigned(31 downto 0);
  signal execute_RS1 : std_logic_vector(31 downto 0);
  attribute keep of execute_RS1 : signal is true;
  attribute syn_keep of execute_RS1 : signal is true;
  signal execute_SHIFT_RIGHT : std_logic_vector(31 downto 0);
  signal zz_decode_RS2_1 : std_logic_vector(31 downto 0);
  signal execute_SHIFT_CTRL : ShiftCtrlEnum_seq_type;
  signal zz_execute_SHIFT_CTRL : ShiftCtrlEnum_seq_type;
  signal execute_SRC_LESS_UNSIGNED : std_logic;
  signal execute_SRC2_FORCE_ZERO : std_logic;
  signal execute_SRC_USE_SUB_LESS : std_logic;
  signal zz_execute_SRC2 : unsigned(31 downto 0);
  signal execute_SRC2_CTRL : Src2CtrlEnum_seq_type;
  signal zz_execute_SRC2_CTRL : Src2CtrlEnum_seq_type;
  signal execute_SRC1_CTRL : Src1CtrlEnum_seq_type;
  signal zz_execute_SRC1_CTRL : Src1CtrlEnum_seq_type;
  signal decode_SRC_USE_SUB_LESS : std_logic;
  signal decode_SRC_ADD_ZERO : std_logic;
  signal execute_SRC_ADD_SUB : std_logic_vector(31 downto 0);
  signal execute_SRC_LESS : std_logic;
  signal execute_ALU_CTRL : AluCtrlEnum_seq_type;
  signal zz_execute_ALU_CTRL : AluCtrlEnum_seq_type;
  signal execute_SRC2 : std_logic_vector(31 downto 0);
  signal execute_SRC1 : std_logic_vector(31 downto 0);
  signal execute_ALU_BITWISE_CTRL : AluBitwiseCtrlEnum_seq_type;
  signal zz_execute_ALU_BITWISE_CTRL : AluBitwiseCtrlEnum_seq_type;
  signal zz_lastStageRegFileWrite_payload_address : std_logic_vector(31 downto 0);
  signal zz_lastStageRegFileWrite_valid : std_logic;
  signal zz_1 : std_logic;
  signal decode_INSTRUCTION_ANTICIPATED : std_logic_vector(31 downto 0);
  signal decode_REGFILE_WRITE_VALID : std_logic;
  signal decode_LEGAL_INSTRUCTION : std_logic;
  signal zz_decode_ENV_CTRL_1 : EnvCtrlEnum_seq_type;
  signal zz_decode_BRANCH_CTRL_1 : BranchCtrlEnum_seq_type;
  signal zz_decode_SHIFT_CTRL_1 : ShiftCtrlEnum_seq_type;
  signal zz_decode_ALU_BITWISE_CTRL_1 : AluBitwiseCtrlEnum_seq_type;
  signal zz_decode_SRC2_CTRL_1 : Src2CtrlEnum_seq_type;
  signal zz_decode_ALU_CTRL_1 : AluCtrlEnum_seq_type;
  signal zz_decode_SRC1_CTRL_1 : Src1CtrlEnum_seq_type;
  signal zz_decode_RS2_2 : std_logic_vector(31 downto 0);
  signal writeBack_MEMORY_WR : std_logic;
  signal writeBack_MEMORY_STORE_DATA_RF : std_logic_vector(31 downto 0);
  signal writeBack_REGFILE_WRITE_DATA : std_logic_vector(31 downto 0);
  signal writeBack_MEMORY_ENABLE : std_logic;
  signal memory_REGFILE_WRITE_DATA : std_logic_vector(31 downto 0);
  signal memory_MEMORY_ENABLE : std_logic;
  signal execute_MEMORY_FORCE_CONSTISTENCY : std_logic;
  signal execute_MEMORY_MANAGMENT : std_logic;
  signal execute_RS2 : std_logic_vector(31 downto 0);
  attribute keep of execute_RS2 : signal is true;
  attribute syn_keep of execute_RS2 : signal is true;
  signal execute_MEMORY_WR : std_logic;
  signal execute_SRC_ADD : std_logic_vector(31 downto 0);
  signal execute_MEMORY_ENABLE : std_logic;
  signal execute_INSTRUCTION : std_logic_vector(31 downto 0);
  signal decode_MEMORY_ENABLE : std_logic;
  signal decode_FLUSH_ALL : std_logic;
  signal IBusCachedPlugin_rsp_issueDetected_4 : std_logic;
  signal IBusCachedPlugin_rsp_issueDetected_3 : std_logic;
  signal IBusCachedPlugin_rsp_issueDetected_2 : std_logic;
  signal IBusCachedPlugin_rsp_issueDetected_1 : std_logic;
  signal decode_INSTRUCTION : std_logic_vector(31 downto 0);
  signal memory_PREDICTION_CONTEXT_hazard : std_logic;
  signal memory_PREDICTION_CONTEXT_hit : std_logic;
  signal memory_PREDICTION_CONTEXT_line_source : std_logic_vector(21 downto 0);
  signal memory_PREDICTION_CONTEXT_line_branchWish : unsigned(1 downto 0);
  signal memory_PREDICTION_CONTEXT_line_target : unsigned(31 downto 0);
  signal zz_2 : std_logic;
  signal zz_memory_to_writeBack_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal decode_PC : unsigned(31 downto 0);
  signal writeBack_PC : unsigned(31 downto 0);
  signal writeBack_INSTRUCTION : std_logic_vector(31 downto 0);
  signal decode_arbitration_haltItself : std_logic;
  signal decode_arbitration_haltByOther : std_logic;
  signal decode_arbitration_removeIt : std_logic;
  signal decode_arbitration_flushIt : std_logic;
  signal decode_arbitration_flushNext : std_logic;
  signal decode_arbitration_isValid : std_logic;
  signal decode_arbitration_isStuck : std_logic;
  signal decode_arbitration_isStuckByOthers : std_logic;
  signal decode_arbitration_isFlushed : std_logic;
  signal decode_arbitration_isMoving : std_logic;
  signal decode_arbitration_isFiring : std_logic;
  signal execute_arbitration_haltItself : std_logic;
  signal execute_arbitration_haltByOther : std_logic;
  signal execute_arbitration_removeIt : std_logic;
  signal execute_arbitration_flushIt : std_logic;
  signal execute_arbitration_flushNext : std_logic;
  signal execute_arbitration_isValid : std_logic;
  signal execute_arbitration_isStuck : std_logic;
  signal execute_arbitration_isStuckByOthers : std_logic;
  signal execute_arbitration_isFlushed : std_logic;
  signal execute_arbitration_isMoving : std_logic;
  signal execute_arbitration_isFiring : std_logic;
  signal memory_arbitration_haltItself : std_logic;
  signal memory_arbitration_haltByOther : std_logic;
  signal memory_arbitration_removeIt : std_logic;
  signal memory_arbitration_flushIt : std_logic;
  signal memory_arbitration_flushNext : std_logic;
  signal memory_arbitration_isValid : std_logic;
  signal memory_arbitration_isStuck : std_logic;
  signal memory_arbitration_isStuckByOthers : std_logic;
  signal memory_arbitration_isFlushed : std_logic;
  signal memory_arbitration_isMoving : std_logic;
  signal memory_arbitration_isFiring : std_logic;
  signal writeBack_arbitration_haltItself : std_logic;
  signal writeBack_arbitration_haltByOther : std_logic;
  signal writeBack_arbitration_removeIt : std_logic;
  signal writeBack_arbitration_flushIt : std_logic;
  signal writeBack_arbitration_flushNext : std_logic;
  signal writeBack_arbitration_isValid : std_logic;
  signal writeBack_arbitration_isStuck : std_logic;
  signal writeBack_arbitration_isStuckByOthers : std_logic;
  signal writeBack_arbitration_isFlushed : std_logic;
  signal writeBack_arbitration_isMoving : std_logic;
  signal writeBack_arbitration_isFiring : std_logic;
  signal lastStageInstruction : std_logic_vector(31 downto 0);
  signal lastStagePc : unsigned(31 downto 0);
  signal lastStageIsValid : std_logic;
  signal lastStageIsFiring : std_logic;
  signal IBusCachedPlugin_fetcherHalt : std_logic;
  signal IBusCachedPlugin_incomingInstruction : std_logic;
  signal IBusCachedPlugin_fetchPrediction_cmd_hadBranch : std_logic;
  signal IBusCachedPlugin_fetchPrediction_cmd_targetPc : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPrediction_rsp_wasRight : std_logic;
  signal IBusCachedPlugin_fetchPrediction_rsp_finalPc : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPrediction_rsp_sourceLastWord : unsigned(31 downto 0);
  signal IBusCachedPlugin_pcValids_0 : std_logic;
  signal IBusCachedPlugin_pcValids_1 : std_logic;
  signal IBusCachedPlugin_pcValids_2 : std_logic;
  signal IBusCachedPlugin_pcValids_3 : std_logic;
  signal IBusCachedPlugin_decodeExceptionPort_valid : std_logic;
  signal IBusCachedPlugin_decodeExceptionPort_payload_code : unsigned(3 downto 0);
  signal IBusCachedPlugin_decodeExceptionPort_payload_badAddr : unsigned(31 downto 0);
  signal IBusCachedPlugin_mmuBus_cmd_0_isValid : std_logic;
  signal IBusCachedPlugin_mmuBus_cmd_0_isStuck : std_logic;
  signal IBusCachedPlugin_mmuBus_cmd_0_virtualAddress : unsigned(31 downto 0);
  signal IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_physicalAddress : unsigned(31 downto 0);
  signal IBusCachedPlugin_mmuBus_rsp_isIoAccess : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_isPaging : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_allowRead : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_allowWrite : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_allowExecute : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_exception : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_refilling : std_logic;
  signal IBusCachedPlugin_mmuBus_rsp_bypassTranslation : std_logic;
  signal IBusCachedPlugin_mmuBus_end : std_logic;
  signal IBusCachedPlugin_mmuBus_busy : std_logic;
  signal DBusCachedPlugin_mmuBus_cmd_0_isValid : std_logic;
  signal DBusCachedPlugin_mmuBus_cmd_0_isStuck : std_logic;
  signal DBusCachedPlugin_mmuBus_cmd_0_virtualAddress : unsigned(31 downto 0);
  signal DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_physicalAddress : unsigned(31 downto 0);
  signal DBusCachedPlugin_mmuBus_rsp_isIoAccess : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_isPaging : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_allowRead : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_allowWrite : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_allowExecute : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_exception : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_refilling : std_logic;
  signal DBusCachedPlugin_mmuBus_rsp_bypassTranslation : std_logic;
  signal DBusCachedPlugin_mmuBus_end : std_logic;
  signal DBusCachedPlugin_mmuBus_busy : std_logic;
  signal DBusCachedPlugin_redoBranch_valid : std_logic;
  signal DBusCachedPlugin_redoBranch_payload : unsigned(31 downto 0);
  signal DBusCachedPlugin_exceptionBus_valid : std_logic;
  signal DBusCachedPlugin_exceptionBus_payload_code : unsigned(3 downto 0);
  signal DBusCachedPlugin_exceptionBus_payload_badAddr : unsigned(31 downto 0);
  signal zz_when_DBusCachedPlugin_l390 : std_logic;
  signal decodeExceptionPort_valid : std_logic;
  signal decodeExceptionPort_payload_code : unsigned(3 downto 0);
  signal decodeExceptionPort_payload_badAddr : unsigned(31 downto 0);
  signal BranchPlugin_jumpInterface_valid : std_logic;
  signal BranchPlugin_jumpInterface_payload : unsigned(31 downto 0);
  signal BranchPlugin_branchExceptionPort_valid : std_logic;
  signal BranchPlugin_branchExceptionPort_payload_code : unsigned(3 downto 0);
  signal BranchPlugin_branchExceptionPort_payload_badAddr : unsigned(31 downto 0);
  signal CsrPlugin_csrMapping_readDataSignal : std_logic_vector(31 downto 0);
  signal CsrPlugin_csrMapping_readDataInit : std_logic_vector(31 downto 0);
  signal CsrPlugin_csrMapping_writeDataSignal : std_logic_vector(31 downto 0);
  signal CsrPlugin_csrMapping_allowCsrSignal : std_logic;
  signal CsrPlugin_csrMapping_hazardFree : std_logic;
  signal CsrPlugin_inWfi : std_logic;
  signal CsrPlugin_thirdPartyWake : std_logic;
  signal CsrPlugin_jumpInterface_valid : std_logic;
  signal CsrPlugin_jumpInterface_payload : unsigned(31 downto 0);
  signal CsrPlugin_exceptionPendings_0 : std_logic;
  signal CsrPlugin_exceptionPendings_1 : std_logic;
  signal CsrPlugin_exceptionPendings_2 : std_logic;
  signal CsrPlugin_exceptionPendings_3 : std_logic;
  signal contextSwitching : std_logic;
  signal CsrPlugin_privilege : unsigned(1 downto 0);
  signal CsrPlugin_forceMachineWire : std_logic;
  signal CsrPlugin_allowInterrupts : std_logic;
  signal CsrPlugin_allowException : std_logic;
  signal CsrPlugin_allowEbreakException : std_logic;
  signal IBusCachedPlugin_injectionPort_valid : std_logic;
  signal IBusCachedPlugin_injectionPort_ready : std_logic;
  signal IBusCachedPlugin_injectionPort_payload : std_logic_vector(31 downto 0);
  signal IBusCachedPlugin_externalFlush : std_logic;
  signal IBusCachedPlugin_jump_pcLoad_valid : std_logic;
  signal IBusCachedPlugin_jump_pcLoad_payload : unsigned(31 downto 0);
  signal zz_IBusCachedPlugin_jump_pcLoad_payload : unsigned(2 downto 0);
  signal zz_IBusCachedPlugin_jump_pcLoad_payload_1 : std_logic_vector(2 downto 0);
  signal zz_IBusCachedPlugin_jump_pcLoad_payload_2 : std_logic;
  signal zz_IBusCachedPlugin_jump_pcLoad_payload_3 : std_logic;
  signal IBusCachedPlugin_fetchPc_output_valid : std_logic;
  signal IBusCachedPlugin_fetchPc_output_ready : std_logic;
  signal IBusCachedPlugin_fetchPc_output_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPc_pcReg : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPc_correction : std_logic;
  signal IBusCachedPlugin_fetchPc_correctionReg : std_logic;
  signal IBusCachedPlugin_fetchPc_output_fire : std_logic;
  signal IBusCachedPlugin_fetchPc_corrected : std_logic;
  signal IBusCachedPlugin_fetchPc_pcRegPropagate : std_logic;
  signal IBusCachedPlugin_fetchPc_booted : std_logic;
  signal IBusCachedPlugin_fetchPc_inc : std_logic;
  signal when_Fetcher_l131 : std_logic;
  signal IBusCachedPlugin_fetchPc_output_fire_1 : std_logic;
  signal when_Fetcher_l131_1 : std_logic;
  signal IBusCachedPlugin_fetchPc_pc : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPc_predictionPcLoad_valid : std_logic;
  signal IBusCachedPlugin_fetchPc_predictionPcLoad_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPc_redo_valid : std_logic;
  signal IBusCachedPlugin_fetchPc_redo_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_fetchPc_flushed : std_logic;
  signal when_Fetcher_l158 : std_logic;
  signal IBusCachedPlugin_iBusRsp_redoFetch : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_input_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_input_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_input_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_0_output_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_output_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_output_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_0_halt : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_input_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_input_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_input_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_1_output_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_output_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_output_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_1_halt : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_2_input_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_2_input_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_2_input_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_2_output_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_2_output_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_2_output_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_2_halt : std_logic;
  signal zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready : std_logic;
  signal zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready : std_logic;
  signal zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_flush : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_payload : unsigned(31 downto 0);
  signal zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid : std_logic;
  signal zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload : unsigned(31 downto 0);
  signal zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid : std_logic;
  signal zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_readyForError : std_logic;
  signal IBusCachedPlugin_iBusRsp_output_valid : std_logic;
  signal IBusCachedPlugin_iBusRsp_output_ready : std_logic;
  signal IBusCachedPlugin_iBusRsp_output_payload_pc : unsigned(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_output_payload_rsp_error : std_logic;
  signal IBusCachedPlugin_iBusRsp_output_payload_rsp_inst : std_logic_vector(31 downto 0);
  signal IBusCachedPlugin_iBusRsp_output_payload_isRvc : std_logic;
  signal when_Fetcher_l240 : std_logic;
  signal when_Fetcher_l320 : std_logic;
  signal IBusCachedPlugin_injector_nextPcCalc_valids_0 : std_logic;
  signal when_Fetcher_l329 : std_logic;
  signal IBusCachedPlugin_injector_nextPcCalc_valids_1 : std_logic;
  signal when_Fetcher_l329_1 : std_logic;
  signal IBusCachedPlugin_injector_nextPcCalc_valids_2 : std_logic;
  signal when_Fetcher_l329_2 : std_logic;
  signal IBusCachedPlugin_injector_nextPcCalc_valids_3 : std_logic;
  signal when_Fetcher_l329_3 : std_logic;
  signal IBusCachedPlugin_injector_nextPcCalc_valids_4 : std_logic;
  signal when_Fetcher_l329_4 : std_logic;
  signal IBusCachedPlugin_predictor_historyWriteDelayPatched_valid : std_logic;
  signal IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_address : unsigned(7 downto 0);
  signal IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_target : unsigned(31 downto 0);
  signal IBusCachedPlugin_predictor_historyWrite_valid : std_logic;
  signal IBusCachedPlugin_predictor_historyWrite_payload_address : unsigned(7 downto 0);
  signal IBusCachedPlugin_predictor_historyWrite_payload_data_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_historyWrite_payload_data_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_historyWrite_payload_data_target : unsigned(31 downto 0);
  signal IBusCachedPlugin_predictor_writeLast_valid : std_logic;
  signal IBusCachedPlugin_predictor_writeLast_payload_address : unsigned(7 downto 0);
  signal IBusCachedPlugin_predictor_writeLast_payload_data_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_writeLast_payload_data_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_writeLast_payload_data_target : unsigned(31 downto 0);
  signal zz_IBusCachedPlugin_predictor_buffer_line_source : unsigned(29 downto 0);
  signal IBusCachedPlugin_predictor_buffer_line_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_buffer_line_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_buffer_line_target : unsigned(31 downto 0);
  signal zz_IBusCachedPlugin_predictor_buffer_line_source_1 : std_logic_vector(55 downto 0);
  signal IBusCachedPlugin_predictor_buffer_pcCorrected : std_logic;
  signal IBusCachedPlugin_predictor_buffer_hazard : std_logic;
  signal IBusCachedPlugin_predictor_line_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_line_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_line_target : unsigned(31 downto 0);
  signal IBusCachedPlugin_predictor_buffer_hazard_regNextWhen : std_logic;
  signal IBusCachedPlugin_predictor_hazard : std_logic;
  signal IBusCachedPlugin_predictor_hit : std_logic;
  signal IBusCachedPlugin_predictor_fetchContext_hazard : std_logic;
  signal IBusCachedPlugin_predictor_fetchContext_hit : std_logic;
  signal IBusCachedPlugin_predictor_fetchContext_line_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_fetchContext_line_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_fetchContext_line_target : unsigned(31 downto 0);
  signal IBusCachedPlugin_predictor_iBusRspContext_hazard : std_logic;
  signal IBusCachedPlugin_predictor_iBusRspContext_hit : std_logic;
  signal IBusCachedPlugin_predictor_iBusRspContext_line_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_iBusRspContext_line_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_iBusRspContext_line_target : unsigned(31 downto 0);
  signal IBusCachedPlugin_predictor_iBusRspContextOutput_hazard : std_logic;
  signal IBusCachedPlugin_predictor_iBusRspContextOutput_hit : std_logic;
  signal IBusCachedPlugin_predictor_iBusRspContextOutput_line_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_iBusRspContextOutput_line_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_iBusRspContextOutput_line_target : unsigned(31 downto 0);
  signal IBusCachedPlugin_predictor_injectorContext_hazard : std_logic;
  signal IBusCachedPlugin_predictor_injectorContext_hit : std_logic;
  signal IBusCachedPlugin_predictor_injectorContext_line_source : std_logic_vector(21 downto 0);
  signal IBusCachedPlugin_predictor_injectorContext_line_branchWish : unsigned(1 downto 0);
  signal IBusCachedPlugin_predictor_injectorContext_line_target : unsigned(31 downto 0);
  signal when_Fetcher_l596 : std_logic;
  signal zz_IBusCachedPlugin_rspCounter : unsigned(31 downto 0);
  signal IBusCachedPlugin_rspCounter : unsigned(31 downto 0);
  signal IBusCachedPlugin_s0_tightlyCoupledHit : std_logic;
  signal IBusCachedPlugin_s1_tightlyCoupledHit : std_logic;
  signal IBusCachedPlugin_s2_tightlyCoupledHit : std_logic;
  signal IBusCachedPlugin_rsp_iBusRspOutputHalt : std_logic;
  signal IBusCachedPlugin_rsp_issueDetected : std_logic;
  signal IBusCachedPlugin_rsp_redoFetch : std_logic;
  signal when_IBusCachedPlugin_l239 : std_logic;
  signal when_IBusCachedPlugin_l244 : std_logic;
  signal when_IBusCachedPlugin_l250 : std_logic;
  signal when_IBusCachedPlugin_l256 : std_logic;
  signal when_IBusCachedPlugin_l267 : std_logic;
  signal zz_DBusCachedPlugin_rspCounter : unsigned(31 downto 0);
  signal DBusCachedPlugin_rspCounter : unsigned(31 downto 0);
  signal when_DBusCachedPlugin_l307 : std_logic;
  signal execute_DBusCachedPlugin_size : unsigned(1 downto 0);
  signal zz_execute_MEMORY_STORE_DATA_RF : std_logic_vector(31 downto 0);
  signal dataCache_1_io_cpu_flush_isStall : std_logic;
  signal when_DBusCachedPlugin_l347 : std_logic;
  signal when_DBusCachedPlugin_l363 : std_logic;
  signal when_DBusCachedPlugin_l390 : std_logic;
  signal when_DBusCachedPlugin_l442 : std_logic;
  signal when_DBusCachedPlugin_l462 : std_logic;
  signal writeBack_DBusCachedPlugin_rspSplits_0 : std_logic_vector(7 downto 0);
  signal writeBack_DBusCachedPlugin_rspSplits_1 : std_logic_vector(7 downto 0);
  signal writeBack_DBusCachedPlugin_rspSplits_2 : std_logic_vector(7 downto 0);
  signal writeBack_DBusCachedPlugin_rspSplits_3 : std_logic_vector(7 downto 0);
  signal writeBack_DBusCachedPlugin_rspShifted : std_logic_vector(31 downto 0);
  signal writeBack_DBusCachedPlugin_rspRf : std_logic_vector(31 downto 0);
  signal switch_Misc_l204 : std_logic_vector(1 downto 0);
  signal zz_writeBack_DBusCachedPlugin_rspFormated : std_logic;
  signal zz_writeBack_DBusCachedPlugin_rspFormated_1 : std_logic_vector(31 downto 0);
  signal zz_writeBack_DBusCachedPlugin_rspFormated_2 : std_logic;
  signal zz_writeBack_DBusCachedPlugin_rspFormated_3 : std_logic_vector(31 downto 0);
  signal writeBack_DBusCachedPlugin_rspFormated : std_logic_vector(31 downto 0);
  signal when_DBusCachedPlugin_l488 : std_logic;
  signal zz_decode_ENV_CTRL_2 : std_logic_vector(31 downto 0);
  signal zz_decode_ENV_CTRL_3 : std_logic;
  signal zz_decode_ENV_CTRL_4 : std_logic;
  signal zz_decode_ENV_CTRL_5 : std_logic;
  signal zz_decode_ENV_CTRL_6 : std_logic;
  signal zz_decode_ENV_CTRL_7 : std_logic;
  signal zz_decode_ENV_CTRL_8 : std_logic;
  signal zz_decode_SRC1_CTRL_2 : Src1CtrlEnum_seq_type;
  signal zz_decode_ALU_CTRL_2 : AluCtrlEnum_seq_type;
  signal zz_decode_SRC2_CTRL_2 : Src2CtrlEnum_seq_type;
  signal zz_decode_ALU_BITWISE_CTRL_2 : AluBitwiseCtrlEnum_seq_type;
  signal zz_decode_SHIFT_CTRL_2 : ShiftCtrlEnum_seq_type;
  signal zz_decode_BRANCH_CTRL_2 : BranchCtrlEnum_seq_type;
  signal zz_decode_ENV_CTRL_9 : EnvCtrlEnum_seq_type;
  signal when_RegFilePlugin_l63 : std_logic;
  signal decode_RegFilePlugin_regFileReadAddress1 : unsigned(4 downto 0);
  signal decode_RegFilePlugin_regFileReadAddress2 : unsigned(4 downto 0);
  signal decode_RegFilePlugin_rs1Data : std_logic_vector(31 downto 0);
  signal decode_RegFilePlugin_rs2Data : std_logic_vector(31 downto 0);
  signal lastStageRegFileWrite_valid : std_logic;
  signal lastStageRegFileWrite_payload_address : unsigned(4 downto 0);
  signal lastStageRegFileWrite_payload_data : std_logic_vector(31 downto 0);
  signal zz_3 : std_logic;
  signal execute_IntAluPlugin_bitwise : std_logic_vector(31 downto 0);
  signal zz_execute_REGFILE_WRITE_DATA : std_logic_vector(31 downto 0);
  signal zz_execute_SRC1 : std_logic_vector(31 downto 0);
  signal zz_execute_SRC2_1 : std_logic;
  signal zz_execute_SRC2_2 : std_logic_vector(19 downto 0);
  signal zz_execute_SRC2_3 : std_logic;
  signal zz_execute_SRC2_4 : std_logic_vector(19 downto 0);
  signal zz_execute_SRC2_5 : std_logic_vector(31 downto 0);
  signal execute_SrcPlugin_addSub : std_logic_vector(31 downto 0);
  signal execute_SrcPlugin_less : std_logic;
  signal execute_FullBarrelShifterPlugin_amplitude : unsigned(4 downto 0);
  signal zz_execute_FullBarrelShifterPlugin_reversed : std_logic_vector(31 downto 0);
  signal execute_FullBarrelShifterPlugin_reversed : std_logic_vector(31 downto 0);
  signal zz_decode_RS2_3 : std_logic_vector(31 downto 0);
  signal execute_MulPlugin_aSigned : std_logic;
  signal execute_MulPlugin_bSigned : std_logic;
  signal execute_MulPlugin_a : std_logic_vector(31 downto 0);
  signal execute_MulPlugin_b : std_logic_vector(31 downto 0);
  signal switch_MulPlugin_l87 : std_logic_vector(1 downto 0);
  signal execute_MulPlugin_aULow : unsigned(15 downto 0);
  signal execute_MulPlugin_bULow : unsigned(15 downto 0);
  signal execute_MulPlugin_aSLow : signed(16 downto 0);
  signal execute_MulPlugin_bSLow : signed(16 downto 0);
  signal execute_MulPlugin_aHigh : signed(16 downto 0);
  signal execute_MulPlugin_bHigh : signed(16 downto 0);
  signal writeBack_MulPlugin_result : signed(65 downto 0);
  signal when_MulPlugin_l147 : std_logic;
  signal switch_MulPlugin_l148 : std_logic_vector(1 downto 0);
  signal memory_DivPlugin_rs1 : unsigned(32 downto 0);
  signal memory_DivPlugin_rs2 : unsigned(31 downto 0);
  signal memory_DivPlugin_accumulator : unsigned(64 downto 0);
  signal memory_DivPlugin_frontendOk : std_logic;
  signal memory_DivPlugin_div_needRevert : std_logic;
  signal memory_DivPlugin_div_counter_willIncrement : std_logic;
  signal memory_DivPlugin_div_counter_willClear : std_logic;
  signal memory_DivPlugin_div_counter_valueNext : unsigned(5 downto 0);
  signal memory_DivPlugin_div_counter_value : unsigned(5 downto 0);
  signal memory_DivPlugin_div_counter_willOverflowIfInc : std_logic;
  signal memory_DivPlugin_div_counter_willOverflow : std_logic;
  signal memory_DivPlugin_div_done : std_logic;
  signal when_MulDivIterativePlugin_l126 : std_logic;
  signal when_MulDivIterativePlugin_l126_1 : std_logic;
  signal memory_DivPlugin_div_result : std_logic_vector(31 downto 0);
  signal when_MulDivIterativePlugin_l128 : std_logic;
  signal when_MulDivIterativePlugin_l129 : std_logic;
  signal when_MulDivIterativePlugin_l132 : std_logic;
  signal zz_memory_DivPlugin_div_stage_0_remainderShifted : unsigned(31 downto 0);
  signal memory_DivPlugin_div_stage_0_remainderShifted : unsigned(32 downto 0);
  signal memory_DivPlugin_div_stage_0_remainderMinusDenominator : unsigned(32 downto 0);
  signal memory_DivPlugin_div_stage_0_outRemainder : unsigned(31 downto 0);
  signal memory_DivPlugin_div_stage_0_outNumerator : unsigned(31 downto 0);
  signal when_MulDivIterativePlugin_l151 : std_logic;
  signal zz_memory_DivPlugin_div_result : unsigned(31 downto 0);
  signal when_MulDivIterativePlugin_l162 : std_logic;
  signal zz_memory_DivPlugin_rs2 : std_logic;
  signal zz_memory_DivPlugin_rs1 : std_logic;
  signal zz_memory_DivPlugin_rs1_1 : std_logic_vector(32 downto 0);
  signal HazardSimplePlugin_src0Hazard : std_logic;
  signal HazardSimplePlugin_src1Hazard : std_logic;
  signal HazardSimplePlugin_writeBackWrites_valid : std_logic;
  signal HazardSimplePlugin_writeBackWrites_payload_address : std_logic_vector(4 downto 0);
  signal HazardSimplePlugin_writeBackWrites_payload_data : std_logic_vector(31 downto 0);
  signal HazardSimplePlugin_writeBackBuffer_valid : std_logic;
  signal HazardSimplePlugin_writeBackBuffer_payload_address : std_logic_vector(4 downto 0);
  signal HazardSimplePlugin_writeBackBuffer_payload_data : std_logic_vector(31 downto 0);
  signal HazardSimplePlugin_addr0Match : std_logic;
  signal HazardSimplePlugin_addr1Match : std_logic;
  signal when_HazardSimplePlugin_l47 : std_logic;
  signal when_HazardSimplePlugin_l48 : std_logic;
  signal when_HazardSimplePlugin_l51 : std_logic;
  signal when_HazardSimplePlugin_l45 : std_logic;
  signal when_HazardSimplePlugin_l57 : std_logic;
  signal when_HazardSimplePlugin_l58 : std_logic;
  signal when_HazardSimplePlugin_l48_1 : std_logic;
  signal when_HazardSimplePlugin_l51_1 : std_logic;
  signal when_HazardSimplePlugin_l45_1 : std_logic;
  signal when_HazardSimplePlugin_l57_1 : std_logic;
  signal when_HazardSimplePlugin_l58_1 : std_logic;
  signal when_HazardSimplePlugin_l48_2 : std_logic;
  signal when_HazardSimplePlugin_l51_2 : std_logic;
  signal when_HazardSimplePlugin_l45_2 : std_logic;
  signal when_HazardSimplePlugin_l57_2 : std_logic;
  signal when_HazardSimplePlugin_l58_2 : std_logic;
  signal when_HazardSimplePlugin_l105 : std_logic;
  signal when_HazardSimplePlugin_l108 : std_logic;
  signal when_HazardSimplePlugin_l113 : std_logic;
  signal execute_BranchPlugin_eq : std_logic;
  signal switch_Misc_l204_1 : std_logic_vector(2 downto 0);
  signal zz_execute_BRANCH_DO : std_logic;
  signal zz_execute_BRANCH_DO_1 : std_logic;
  signal execute_BranchPlugin_branch_src1 : unsigned(31 downto 0);
  signal zz_execute_BRANCH_SRC22 : std_logic;
  signal zz_execute_BRANCH_SRC22_1 : std_logic_vector(10 downto 0);
  signal zz_execute_BRANCH_SRC22_2 : std_logic;
  signal zz_execute_BRANCH_SRC22_3 : std_logic_vector(19 downto 0);
  signal zz_execute_BRANCH_SRC22_4 : std_logic;
  signal zz_execute_BRANCH_SRC22_5 : std_logic_vector(18 downto 0);
  signal zz_execute_BRANCH_SRC22_6 : std_logic_vector(31 downto 0);
  signal execute_BranchPlugin_branchAdder : unsigned(31 downto 0);
  signal memory_BranchPlugin_predictionMissmatch : std_logic;
  signal CsrPlugin_misa_base : unsigned(1 downto 0);
  signal CsrPlugin_misa_extensions : std_logic_vector(25 downto 0);
  signal CsrPlugin_mtvec_mode : std_logic_vector(1 downto 0);
  signal CsrPlugin_mtvec_base : unsigned(29 downto 0);
  signal CsrPlugin_mepc : unsigned(31 downto 0);
  signal CsrPlugin_mstatus_MIE : std_logic;
  signal CsrPlugin_mstatus_MPIE : std_logic;
  signal CsrPlugin_mstatus_MPP : unsigned(1 downto 0);
  signal CsrPlugin_mip_MEIP : std_logic;
  signal CsrPlugin_mip_MTIP : std_logic;
  signal CsrPlugin_mip_MSIP : std_logic;
  signal CsrPlugin_mie_MEIE : std_logic;
  signal CsrPlugin_mie_MTIE : std_logic;
  signal CsrPlugin_mie_MSIE : std_logic;
  signal CsrPlugin_mcause_interrupt : std_logic;
  signal CsrPlugin_mcause_exceptionCode : unsigned(3 downto 0);
  signal CsrPlugin_mtval : unsigned(31 downto 0);
  signal CsrPlugin_mcycle : unsigned(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000";
  signal CsrPlugin_minstret : unsigned(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000";
  signal zz_when_CsrPlugin_l952 : std_logic;
  signal zz_when_CsrPlugin_l952_1 : std_logic;
  signal zz_when_CsrPlugin_l952_2 : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValids_decode : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValids_execute : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValids_memory : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack : std_logic;
  signal CsrPlugin_exceptionPortCtrl_exceptionContext_code : unsigned(3 downto 0);
  signal CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr : unsigned(31 downto 0);
  signal CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped : unsigned(1 downto 0);
  signal CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege : unsigned(1 downto 0);
  signal zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code : unsigned(1 downto 0);
  signal zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 : std_logic;
  signal when_CsrPlugin_l909 : std_logic;
  signal when_CsrPlugin_l909_1 : std_logic;
  signal when_CsrPlugin_l909_2 : std_logic;
  signal when_CsrPlugin_l909_3 : std_logic;
  signal when_CsrPlugin_l922 : std_logic;
  signal CsrPlugin_interrupt_valid : std_logic;
  signal CsrPlugin_interrupt_code : unsigned(3 downto 0);
  signal CsrPlugin_interrupt_targetPrivilege : unsigned(1 downto 0);
  signal when_CsrPlugin_l946 : std_logic;
  signal when_CsrPlugin_l952 : std_logic;
  signal when_CsrPlugin_l952_1 : std_logic;
  signal when_CsrPlugin_l952_2 : std_logic;
  signal CsrPlugin_exception : std_logic;
  signal CsrPlugin_lastStageWasWfi : std_logic;
  signal CsrPlugin_pipelineLiberator_pcValids_0 : std_logic;
  signal CsrPlugin_pipelineLiberator_pcValids_1 : std_logic;
  signal CsrPlugin_pipelineLiberator_pcValids_2 : std_logic;
  signal CsrPlugin_pipelineLiberator_active : std_logic;
  signal when_CsrPlugin_l980 : std_logic;
  signal when_CsrPlugin_l980_1 : std_logic;
  signal when_CsrPlugin_l980_2 : std_logic;
  signal when_CsrPlugin_l985 : std_logic;
  signal CsrPlugin_pipelineLiberator_done : std_logic;
  signal when_CsrPlugin_l991 : std_logic;
  signal CsrPlugin_interruptJump : std_logic;
  signal CsrPlugin_hadException : std_logic;
  signal CsrPlugin_targetPrivilege : unsigned(1 downto 0);
  signal CsrPlugin_trapCause : unsigned(3 downto 0);
  signal CsrPlugin_xtvec_mode : std_logic_vector(1 downto 0);
  signal CsrPlugin_xtvec_base : unsigned(29 downto 0);
  signal when_CsrPlugin_l1019 : std_logic;
  signal when_CsrPlugin_l1064 : std_logic;
  signal switch_CsrPlugin_l1068 : std_logic_vector(1 downto 0);
  signal execute_CsrPlugin_wfiWake : std_logic;
  signal when_CsrPlugin_l1116 : std_logic;
  signal execute_CsrPlugin_blockedBySideEffects : std_logic;
  signal execute_CsrPlugin_illegalAccess : std_logic;
  signal execute_CsrPlugin_illegalInstruction : std_logic;
  signal when_CsrPlugin_l1136 : std_logic;
  signal when_CsrPlugin_l1137 : std_logic;
  signal execute_CsrPlugin_writeInstruction : std_logic;
  signal execute_CsrPlugin_readInstruction : std_logic;
  signal execute_CsrPlugin_writeEnable : std_logic;
  signal execute_CsrPlugin_readEnable : std_logic;
  signal execute_CsrPlugin_readToWriteData : std_logic_vector(31 downto 0);
  signal switch_Misc_l204_2 : std_logic;
  signal zz_CsrPlugin_csrMapping_writeDataSignal : std_logic_vector(31 downto 0);
  signal when_CsrPlugin_l1176 : std_logic;
  signal when_CsrPlugin_l1180 : std_logic;
  signal execute_CsrPlugin_csrAddress : std_logic_vector(11 downto 0);
  signal DebugPlugin_firstCycle : std_logic;
  signal DebugPlugin_secondCycle : std_logic;
  signal DebugPlugin_resetIt : std_logic;
  signal DebugPlugin_haltIt : std_logic;
  signal DebugPlugin_stepIt : std_logic;
  signal DebugPlugin_isPipBusy : std_logic;
  signal DebugPlugin_godmode : std_logic;
  signal when_DebugPlugin_l225 : std_logic;
  signal DebugPlugin_haltedByBreak : std_logic;
  signal DebugPlugin_debugUsed : std_logic;
  signal DebugPlugin_disableEbreak : std_logic;
  signal DebugPlugin_allowEBreak : std_logic;
  signal DebugPlugin_busReadDataReg : std_logic_vector(31 downto 0);
  signal zz_when_DebugPlugin_l244 : std_logic;
  signal when_DebugPlugin_l244 : std_logic;
  signal switch_DebugPlugin_l267 : unsigned(5 downto 0);
  signal when_DebugPlugin_l271 : std_logic;
  signal when_DebugPlugin_l271_1 : std_logic;
  signal when_DebugPlugin_l272 : std_logic;
  signal when_DebugPlugin_l272_1 : std_logic;
  signal when_DebugPlugin_l273 : std_logic;
  signal when_DebugPlugin_l274 : std_logic;
  signal when_DebugPlugin_l275 : std_logic;
  signal when_DebugPlugin_l275_1 : std_logic;
  signal when_DebugPlugin_l295 : std_logic;
  signal when_DebugPlugin_l298 : std_logic;
  signal when_DebugPlugin_l311 : std_logic;
  signal DebugPlugin_resetIt_regNext : std_logic;
  signal when_DebugPlugin_l327 : std_logic;
  signal when_Pipeline_l124 : std_logic;
  signal decode_to_execute_PC : unsigned(31 downto 0);
  signal when_Pipeline_l124_1 : std_logic;
  signal execute_to_memory_PC : unsigned(31 downto 0);
  signal when_Pipeline_l124_2 : std_logic;
  signal memory_to_writeBack_PC : unsigned(31 downto 0);
  signal when_Pipeline_l124_3 : std_logic;
  signal decode_to_execute_INSTRUCTION : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_4 : std_logic;
  signal execute_to_memory_INSTRUCTION : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_5 : std_logic;
  signal memory_to_writeBack_INSTRUCTION : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_6 : std_logic;
  signal decode_to_execute_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal when_Pipeline_l124_7 : std_logic;
  signal execute_to_memory_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal when_Pipeline_l124_8 : std_logic;
  signal memory_to_writeBack_FORMAL_PC_NEXT : unsigned(31 downto 0);
  signal when_Pipeline_l124_9 : std_logic;
  signal decode_to_execute_PREDICTION_CONTEXT_hazard : std_logic;
  signal decode_to_execute_PREDICTION_CONTEXT_hit : std_logic;
  signal decode_to_execute_PREDICTION_CONTEXT_line_source : std_logic_vector(21 downto 0);
  signal decode_to_execute_PREDICTION_CONTEXT_line_branchWish : unsigned(1 downto 0);
  signal decode_to_execute_PREDICTION_CONTEXT_line_target : unsigned(31 downto 0);
  signal when_Pipeline_l124_10 : std_logic;
  signal execute_to_memory_PREDICTION_CONTEXT_hazard : std_logic;
  signal execute_to_memory_PREDICTION_CONTEXT_hit : std_logic;
  signal execute_to_memory_PREDICTION_CONTEXT_line_source : std_logic_vector(21 downto 0);
  signal execute_to_memory_PREDICTION_CONTEXT_line_branchWish : unsigned(1 downto 0);
  signal execute_to_memory_PREDICTION_CONTEXT_line_target : unsigned(31 downto 0);
  signal when_Pipeline_l124_11 : std_logic;
  signal decode_to_execute_MEMORY_FORCE_CONSTISTENCY : std_logic;
  signal when_Pipeline_l124_12 : std_logic;
  signal decode_to_execute_SRC1_CTRL : Src1CtrlEnum_seq_type;
  signal when_Pipeline_l124_13 : std_logic;
  signal decode_to_execute_SRC_USE_SUB_LESS : std_logic;
  signal when_Pipeline_l124_14 : std_logic;
  signal decode_to_execute_MEMORY_ENABLE : std_logic;
  signal when_Pipeline_l124_15 : std_logic;
  signal execute_to_memory_MEMORY_ENABLE : std_logic;
  signal when_Pipeline_l124_16 : std_logic;
  signal memory_to_writeBack_MEMORY_ENABLE : std_logic;
  signal when_Pipeline_l124_17 : std_logic;
  signal decode_to_execute_ALU_CTRL : AluCtrlEnum_seq_type;
  signal when_Pipeline_l124_18 : std_logic;
  signal decode_to_execute_SRC2_CTRL : Src2CtrlEnum_seq_type;
  signal when_Pipeline_l124_19 : std_logic;
  signal decode_to_execute_REGFILE_WRITE_VALID : std_logic;
  signal when_Pipeline_l124_20 : std_logic;
  signal execute_to_memory_REGFILE_WRITE_VALID : std_logic;
  signal when_Pipeline_l124_21 : std_logic;
  signal memory_to_writeBack_REGFILE_WRITE_VALID : std_logic;
  signal when_Pipeline_l124_22 : std_logic;
  signal decode_to_execute_BYPASSABLE_EXECUTE_STAGE : std_logic;
  signal when_Pipeline_l124_23 : std_logic;
  signal decode_to_execute_BYPASSABLE_MEMORY_STAGE : std_logic;
  signal when_Pipeline_l124_24 : std_logic;
  signal execute_to_memory_BYPASSABLE_MEMORY_STAGE : std_logic;
  signal when_Pipeline_l124_25 : std_logic;
  signal decode_to_execute_MEMORY_WR : std_logic;
  signal when_Pipeline_l124_26 : std_logic;
  signal execute_to_memory_MEMORY_WR : std_logic;
  signal when_Pipeline_l124_27 : std_logic;
  signal memory_to_writeBack_MEMORY_WR : std_logic;
  signal when_Pipeline_l124_28 : std_logic;
  signal decode_to_execute_MEMORY_MANAGMENT : std_logic;
  signal when_Pipeline_l124_29 : std_logic;
  signal decode_to_execute_SRC_LESS_UNSIGNED : std_logic;
  signal when_Pipeline_l124_30 : std_logic;
  signal decode_to_execute_ALU_BITWISE_CTRL : AluBitwiseCtrlEnum_seq_type;
  signal when_Pipeline_l124_31 : std_logic;
  signal decode_to_execute_SHIFT_CTRL : ShiftCtrlEnum_seq_type;
  signal when_Pipeline_l124_32 : std_logic;
  signal decode_to_execute_IS_MUL : std_logic;
  signal when_Pipeline_l124_33 : std_logic;
  signal execute_to_memory_IS_MUL : std_logic;
  signal when_Pipeline_l124_34 : std_logic;
  signal memory_to_writeBack_IS_MUL : std_logic;
  signal when_Pipeline_l124_35 : std_logic;
  signal decode_to_execute_IS_DIV : std_logic;
  signal when_Pipeline_l124_36 : std_logic;
  signal execute_to_memory_IS_DIV : std_logic;
  signal when_Pipeline_l124_37 : std_logic;
  signal decode_to_execute_IS_RS1_SIGNED : std_logic;
  signal when_Pipeline_l124_38 : std_logic;
  signal decode_to_execute_IS_RS2_SIGNED : std_logic;
  signal when_Pipeline_l124_39 : std_logic;
  signal decode_to_execute_BRANCH_CTRL : BranchCtrlEnum_seq_type;
  signal when_Pipeline_l124_40 : std_logic;
  signal decode_to_execute_IS_CSR : std_logic;
  signal when_Pipeline_l124_41 : std_logic;
  signal decode_to_execute_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal when_Pipeline_l124_42 : std_logic;
  signal execute_to_memory_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal when_Pipeline_l124_43 : std_logic;
  signal memory_to_writeBack_ENV_CTRL : EnvCtrlEnum_seq_type;
  signal when_Pipeline_l124_44 : std_logic;
  signal decode_to_execute_RS1 : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_45 : std_logic;
  signal decode_to_execute_RS2 : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_46 : std_logic;
  signal decode_to_execute_SRC2_FORCE_ZERO : std_logic;
  signal when_Pipeline_l124_47 : std_logic;
  signal decode_to_execute_CSR_WRITE_OPCODE : std_logic;
  signal when_Pipeline_l124_48 : std_logic;
  signal decode_to_execute_CSR_READ_OPCODE : std_logic;
  signal when_Pipeline_l124_49 : std_logic;
  signal decode_to_execute_DO_EBREAK : std_logic;
  signal when_Pipeline_l124_50 : std_logic;
  signal execute_to_memory_MEMORY_STORE_DATA_RF : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_51 : std_logic;
  signal memory_to_writeBack_MEMORY_STORE_DATA_RF : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_52 : std_logic;
  signal execute_to_memory_REGFILE_WRITE_DATA : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_53 : std_logic;
  signal memory_to_writeBack_REGFILE_WRITE_DATA : std_logic_vector(31 downto 0);
  signal when_Pipeline_l124_54 : std_logic;
  signal execute_to_memory_MUL_LL : unsigned(31 downto 0);
  signal when_Pipeline_l124_55 : std_logic;
  signal execute_to_memory_MUL_LH : signed(33 downto 0);
  signal when_Pipeline_l124_56 : std_logic;
  signal execute_to_memory_MUL_HL : signed(33 downto 0);
  signal when_Pipeline_l124_57 : std_logic;
  signal execute_to_memory_MUL_HH : signed(33 downto 0);
  signal when_Pipeline_l124_58 : std_logic;
  signal memory_to_writeBack_MUL_HH : signed(33 downto 0);
  signal when_Pipeline_l124_59 : std_logic;
  signal execute_to_memory_BRANCH_DO : std_logic;
  signal when_Pipeline_l124_60 : std_logic;
  signal execute_to_memory_BRANCH_CALC : unsigned(31 downto 0);
  signal when_Pipeline_l124_61 : std_logic;
  signal execute_to_memory_NEXT_PC2 : unsigned(31 downto 0);
  signal when_Pipeline_l124_62 : std_logic;
  signal execute_to_memory_TARGET_MISSMATCH2 : std_logic;
  signal when_Pipeline_l124_63 : std_logic;
  signal memory_to_writeBack_MUL_LOW : signed(51 downto 0);
  signal when_Pipeline_l151 : std_logic;
  signal when_Pipeline_l154 : std_logic;
  signal when_Pipeline_l151_1 : std_logic;
  signal when_Pipeline_l154_1 : std_logic;
  signal when_Pipeline_l151_2 : std_logic;
  signal when_Pipeline_l154_2 : std_logic;
  signal switch_Fetcher_l362 : unsigned(2 downto 0);
  signal when_Fetcher_l378 : std_logic;
  signal when_CsrPlugin_l1264 : std_logic;
  signal execute_CsrPlugin_csr_768 : std_logic;
  signal when_CsrPlugin_l1264_1 : std_logic;
  signal execute_CsrPlugin_csr_836 : std_logic;
  signal when_CsrPlugin_l1264_2 : std_logic;
  signal execute_CsrPlugin_csr_772 : std_logic;
  signal when_CsrPlugin_l1264_3 : std_logic;
  signal execute_CsrPlugin_csr_833 : std_logic;
  signal when_CsrPlugin_l1264_4 : std_logic;
  signal execute_CsrPlugin_csr_834 : std_logic;
  signal when_CsrPlugin_l1264_5 : std_logic;
  signal execute_CsrPlugin_csr_835 : std_logic;
  signal zz_CsrPlugin_csrMapping_readDataInit : std_logic_vector(31 downto 0);
  signal zz_CsrPlugin_csrMapping_readDataInit_1 : std_logic_vector(31 downto 0);
  signal zz_CsrPlugin_csrMapping_readDataInit_2 : std_logic_vector(31 downto 0);
  signal zz_CsrPlugin_csrMapping_readDataInit_3 : std_logic_vector(31 downto 0);
  signal zz_CsrPlugin_csrMapping_readDataInit_4 : std_logic_vector(31 downto 0);
  signal zz_CsrPlugin_csrMapping_readDataInit_5 : std_logic_vector(31 downto 0);
  signal when_CsrPlugin_l1297 : std_logic;
  signal when_CsrPlugin_l1302 : std_logic;
  type IBusCachedPlugin_predictor_history_type is array (0 to 255) of std_logic_vector(55 downto 0);
  signal IBusCachedPlugin_predictor_history : IBusCachedPlugin_predictor_history_type;
  type RegFilePlugin_regFile_type is array (0 to 31) of std_logic_vector(31 downto 0);
  signal RegFilePlugin_regFile : RegFilePlugin_regFile_type;
begin
  debug_bus_cmd_ready <= debug_bus_cmd_ready_read_buffer;
  zz_when <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(decodeExceptionPort_valid),pkg_toStdLogicVector(IBusCachedPlugin_decodeExceptionPort_valid)) /= pkg_stdLogicVector("00"));
  zz_IBusCachedPlugin_predictor_history_port <= pkg_cat(std_logic_vector(IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_target),pkg_cat(std_logic_vector(IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_branchWish),IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_source));
  zz_zz_IBusCachedPlugin_predictor_buffer_line_source_1 <= pkg_resize(zz_IBusCachedPlugin_predictor_buffer_line_source,8);
  zz_decode_RegFilePlugin_rs1Data <= pkg_toStdLogic(true);
  zz_decode_RegFilePlugin_rs2Data <= pkg_toStdLogic(true);
  zz_IBusCachedPlugin_jump_pcLoad_payload_5 <= unsigned(pkg_cat(pkg_toStdLogicVector(zz_IBusCachedPlugin_jump_pcLoad_payload_3),pkg_toStdLogicVector(zz_IBusCachedPlugin_jump_pcLoad_payload_2)));
  zz_writeBack_DBusCachedPlugin_rspShifted_1 <= pkg_extract(dataCache_1_io_cpu_writeBack_address,1,0);
  zz_writeBack_DBusCachedPlugin_rspShifted_3 <= pkg_extract(dataCache_1_io_cpu_writeBack_address,1,1);
  zz_decode_LEGAL_INSTRUCTION <= pkg_stdLogicVector("00000000000000000001000001101111");
  zz_decode_LEGAL_INSTRUCTION_1 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000001000001111111"));
  zz_decode_LEGAL_INSTRUCTION_2 <= pkg_stdLogicVector("00000000000000000001000001110011");
  zz_decode_LEGAL_INSTRUCTION_3 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000010000001111111")) = pkg_stdLogicVector("00000000000000000010000001110011"));
  zz_decode_LEGAL_INSTRUCTION_4 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000100000001111111")) = pkg_stdLogicVector("00000000000000000100000001100011")));
  zz_decode_LEGAL_INSTRUCTION_5 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000010000001111111")) = pkg_stdLogicVector("00000000000000000010000000010011"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000110000000111111")) = pkg_stdLogicVector("00000000000000000000000000100011"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_decode_LEGAL_INSTRUCTION_6) = pkg_stdLogicVector("00000000000000000000000000000011"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_decode_LEGAL_INSTRUCTION_7 = zz_decode_LEGAL_INSTRUCTION_8)),pkg_cat(pkg_toStdLogicVector(zz_decode_LEGAL_INSTRUCTION_9),pkg_cat(zz_decode_LEGAL_INSTRUCTION_10,zz_decode_LEGAL_INSTRUCTION_11))))));
  zz_decode_LEGAL_INSTRUCTION_6 <= pkg_stdLogicVector("00000000000000000010000001111111");
  zz_decode_LEGAL_INSTRUCTION_7 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000101000001011111"));
  zz_decode_LEGAL_INSTRUCTION_8 <= pkg_stdLogicVector("00000000000000000000000000000011");
  zz_decode_LEGAL_INSTRUCTION_9 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000111000001111011")) = pkg_stdLogicVector("00000000000000000000000001100011"));
  zz_decode_LEGAL_INSTRUCTION_10 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000110000001111111")) = pkg_stdLogicVector("00000000000000000000000000001111")));
  zz_decode_LEGAL_INSTRUCTION_11 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("11111100000000000000000001111111")) = pkg_stdLogicVector("00000000000000000000000000110011"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000001111100000111000001111111")) = pkg_stdLogicVector("00000000000000000101000000001111"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_decode_LEGAL_INSTRUCTION_12) = pkg_stdLogicVector("00000000000000000101000000010011"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_decode_LEGAL_INSTRUCTION_13 = zz_decode_LEGAL_INSTRUCTION_14)),pkg_cat(pkg_toStdLogicVector(zz_decode_LEGAL_INSTRUCTION_15),pkg_cat(zz_decode_LEGAL_INSTRUCTION_16,zz_decode_LEGAL_INSTRUCTION_17))))));
  zz_decode_LEGAL_INSTRUCTION_12 <= pkg_stdLogicVector("10111100000000000111000001111111");
  zz_decode_LEGAL_INSTRUCTION_13 <= (decode_INSTRUCTION and pkg_stdLogicVector("11111100000000000011000001111111"));
  zz_decode_LEGAL_INSTRUCTION_14 <= pkg_stdLogicVector("00000000000000000001000000010011");
  zz_decode_LEGAL_INSTRUCTION_15 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("10111110000000000111000001111111")) = pkg_stdLogicVector("00000000000000000101000000110011"));
  zz_decode_LEGAL_INSTRUCTION_16 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("10111110000000000111000001111111")) = pkg_stdLogicVector("00000000000000000000000000110011")));
  zz_decode_LEGAL_INSTRUCTION_17 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("11011111111111111111111111111111")) = pkg_stdLogicVector("00010000001000000000000001110011"))),pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("11111111111111111111111111111111")) = pkg_stdLogicVector("00000000000100000000000001110011"))));
  zz_zz_decode_ENV_CTRL_2 <= pkg_stdLogicVector("00010000000000000011000001010000");
  zz_zz_decode_ENV_CTRL_2_1 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000100000011000001010000"));
  zz_zz_decode_ENV_CTRL_2_2 <= pkg_stdLogicVector("00000000000000000000000001010000");
  zz_zz_decode_ENV_CTRL_2_3 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_4) = pkg_stdLogicVector("00000000000000000001000001010000")));
  zz_zz_decode_ENV_CTRL_2_5 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_6) = pkg_stdLogicVector("00000000000000000010000001010000")));
  zz_zz_decode_ENV_CTRL_2_7 <= pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_6),pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_8 = zz_zz_decode_ENV_CTRL_2_9)));
  zz_zz_decode_ENV_CTRL_2_10 <= pkg_stdLogicVector("00");
  zz_zz_decode_ENV_CTRL_2_11 <= pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_12 = zz_zz_decode_ENV_CTRL_2_13)) /= pkg_stdLogicVector("0"));
  zz_zz_decode_ENV_CTRL_2_14 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_toStdLogicVector(zz_decode_ENV_CTRL_8) /= pkg_stdLogicVector("0")));
  zz_zz_decode_ENV_CTRL_2_15 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_16 /= zz_zz_decode_ENV_CTRL_2_17)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_18),pkg_cat(zz_zz_decode_ENV_CTRL_2_19,zz_zz_decode_ENV_CTRL_2_21)));
  zz_zz_decode_ENV_CTRL_2_4 <= pkg_stdLogicVector("00000000000000000001000001010000");
  zz_zz_decode_ENV_CTRL_2_6 <= pkg_stdLogicVector("00000000000000000010000001010000");
  zz_zz_decode_ENV_CTRL_2_8 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000011100"));
  zz_zz_decode_ENV_CTRL_2_9 <= pkg_stdLogicVector("00000000000000000000000000000100");
  zz_zz_decode_ENV_CTRL_2_12 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001011000"));
  zz_zz_decode_ENV_CTRL_2_13 <= pkg_stdLogicVector("00000000000000000000000001000000");
  zz_zz_decode_ENV_CTRL_2_16 <= pkg_toStdLogicVector(zz_decode_ENV_CTRL_8);
  zz_zz_decode_ENV_CTRL_2_17 <= pkg_stdLogicVector("0");
  zz_zz_decode_ENV_CTRL_2_18 <= pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000010000000000100000001100100")) = pkg_stdLogicVector("00000010000000000100000000100000"))) /= pkg_stdLogicVector("0"));
  zz_zz_decode_ENV_CTRL_2_19 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_20) = pkg_stdLogicVector("00000010000000000000000000110000"))) /= pkg_stdLogicVector("0")));
  zz_zz_decode_ENV_CTRL_2_21 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_22),pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_23)) /= pkg_stdLogicVector("00"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_24,zz_zz_decode_ENV_CTRL_2_26) /= pkg_stdLogicVector("000"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_31 /= zz_zz_decode_ENV_CTRL_2_33)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_34),pkg_cat(zz_zz_decode_ENV_CTRL_2_37,zz_zz_decode_ENV_CTRL_2_39)))));
  zz_zz_decode_ENV_CTRL_2_20 <= pkg_stdLogicVector("00000010000000000100000001110100");
  zz_zz_decode_ENV_CTRL_2_22 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000111000000110100")) = pkg_stdLogicVector("00000000000000000101000000010000"));
  zz_zz_decode_ENV_CTRL_2_23 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000010000000000111000001100100")) = pkg_stdLogicVector("00000000000000000101000000100000"));
  zz_zz_decode_ENV_CTRL_2_24 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_25) = pkg_stdLogicVector("01000000000000000001000000010000")));
  zz_zz_decode_ENV_CTRL_2_26 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_27 = zz_zz_decode_ENV_CTRL_2_28)),pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_29 = zz_zz_decode_ENV_CTRL_2_30)));
  zz_zz_decode_ENV_CTRL_2_31 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_32) = pkg_stdLogicVector("00000000000000000000000000100100")));
  zz_zz_decode_ENV_CTRL_2_33 <= pkg_stdLogicVector("0");
  zz_zz_decode_ENV_CTRL_2_34 <= pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_35 = zz_zz_decode_ENV_CTRL_2_36)) /= pkg_stdLogicVector("0"));
  zz_zz_decode_ENV_CTRL_2_37 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_38) /= pkg_stdLogicVector("0")));
  zz_zz_decode_ENV_CTRL_2_39 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_40 /= zz_zz_decode_ENV_CTRL_2_45)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_46),pkg_cat(zz_zz_decode_ENV_CTRL_2_49,zz_zz_decode_ENV_CTRL_2_54)));
  zz_zz_decode_ENV_CTRL_2_25 <= pkg_stdLogicVector("01000000000000000011000001010100");
  zz_zz_decode_ENV_CTRL_2_27 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000111000000110100"));
  zz_zz_decode_ENV_CTRL_2_28 <= pkg_stdLogicVector("00000000000000000001000000010000");
  zz_zz_decode_ENV_CTRL_2_29 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000010000000000111000001010100"));
  zz_zz_decode_ENV_CTRL_2_30 <= pkg_stdLogicVector("00000000000000000001000000010000");
  zz_zz_decode_ENV_CTRL_2_32 <= pkg_stdLogicVector("00000000000000000000000001100100");
  zz_zz_decode_ENV_CTRL_2_35 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000001000000000000"));
  zz_zz_decode_ENV_CTRL_2_36 <= pkg_stdLogicVector("00000000000000000001000000000000");
  zz_zz_decode_ENV_CTRL_2_38 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000011000000000000")) = pkg_stdLogicVector("00000000000000000010000000000000"));
  zz_zz_decode_ENV_CTRL_2_40 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_41 = zz_zz_decode_ENV_CTRL_2_42)),pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_43 = zz_zz_decode_ENV_CTRL_2_44)));
  zz_zz_decode_ENV_CTRL_2_45 <= pkg_stdLogicVector("00");
  zz_zz_decode_ENV_CTRL_2_46 <= pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_47 = zz_zz_decode_ENV_CTRL_2_48)) /= pkg_stdLogicVector("0"));
  zz_zz_decode_ENV_CTRL_2_49 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_50,zz_zz_decode_ENV_CTRL_2_52) /= pkg_stdLogicVector("00")));
  zz_zz_decode_ENV_CTRL_2_54 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_55 /= zz_zz_decode_ENV_CTRL_2_59)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_60),pkg_cat(zz_zz_decode_ENV_CTRL_2_63,zz_zz_decode_ENV_CTRL_2_73)));
  zz_zz_decode_ENV_CTRL_2_41 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000010000000010000"));
  zz_zz_decode_ENV_CTRL_2_42 <= pkg_stdLogicVector("00000000000000000010000000000000");
  zz_zz_decode_ENV_CTRL_2_43 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000101000000000000"));
  zz_zz_decode_ENV_CTRL_2_44 <= pkg_stdLogicVector("00000000000000000001000000000000");
  zz_zz_decode_ENV_CTRL_2_47 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000100000001001000"));
  zz_zz_decode_ENV_CTRL_2_48 <= pkg_stdLogicVector("00000000000000000100000000001000");
  zz_zz_decode_ENV_CTRL_2_50 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_51) = pkg_stdLogicVector("00000000000000000000000000100000")));
  zz_zz_decode_ENV_CTRL_2_52 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_53) = pkg_stdLogicVector("00000000000000000000000000100000")));
  zz_zz_decode_ENV_CTRL_2_55 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_56 = zz_zz_decode_ENV_CTRL_2_57)),pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_4),pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_58)));
  zz_zz_decode_ENV_CTRL_2_59 <= pkg_stdLogicVector("000");
  zz_zz_decode_ENV_CTRL_2_60 <= pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_61 = zz_zz_decode_ENV_CTRL_2_62)) /= pkg_stdLogicVector("0"));
  zz_zz_decode_ENV_CTRL_2_63 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_64,zz_zz_decode_ENV_CTRL_2_66) /= pkg_stdLogicVector("00000")));
  zz_zz_decode_ENV_CTRL_2_73 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_74 /= zz_zz_decode_ENV_CTRL_2_77)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_78),pkg_cat(zz_zz_decode_ENV_CTRL_2_91,zz_zz_decode_ENV_CTRL_2_96)));
  zz_zz_decode_ENV_CTRL_2_51 <= pkg_stdLogicVector("00000000000000000000000000110100");
  zz_zz_decode_ENV_CTRL_2_53 <= pkg_stdLogicVector("00000000000000000000000001100100");
  zz_zz_decode_ENV_CTRL_2_56 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001010000"));
  zz_zz_decode_ENV_CTRL_2_57 <= pkg_stdLogicVector("00000000000000000000000001000000");
  zz_zz_decode_ENV_CTRL_2_58 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000100000011000001000000")) = pkg_stdLogicVector("00000000000000000000000001000000"));
  zz_zz_decode_ENV_CTRL_2_61 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000100000"));
  zz_zz_decode_ENV_CTRL_2_62 <= pkg_stdLogicVector("00000000000000000000000000100000");
  zz_zz_decode_ENV_CTRL_2_64 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_65) = pkg_stdLogicVector("00000000000000000000000001000000")));
  zz_zz_decode_ENV_CTRL_2_66 <= pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_5),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_67),pkg_cat(zz_zz_decode_ENV_CTRL_2_69,zz_zz_decode_ENV_CTRL_2_70)));
  zz_zz_decode_ENV_CTRL_2_74 <= pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_5),pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_7),pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_75)));
  zz_zz_decode_ENV_CTRL_2_77 <= pkg_stdLogicVector("000");
  zz_zz_decode_ENV_CTRL_2_78 <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_6),pkg_cat(zz_zz_decode_ENV_CTRL_2_79,zz_zz_decode_ENV_CTRL_2_82)) /= pkg_stdLogicVector("000000"));
  zz_zz_decode_ENV_CTRL_2_91 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_92,zz_zz_decode_ENV_CTRL_2_93) /= pkg_stdLogicVector("00")));
  zz_zz_decode_ENV_CTRL_2_96 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_97 /= zz_zz_decode_ENV_CTRL_2_100)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_101),pkg_cat(zz_zz_decode_ENV_CTRL_2_104,zz_zz_decode_ENV_CTRL_2_109)));
  zz_zz_decode_ENV_CTRL_2_65 <= pkg_stdLogicVector("00000000000000000000000001000000");
  zz_zz_decode_ENV_CTRL_2_67 <= pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_68) = pkg_stdLogicVector("00000000000000000100000000100000"));
  zz_zz_decode_ENV_CTRL_2_69 <= pkg_toStdLogicVector(zz_decode_ENV_CTRL_7);
  zz_zz_decode_ENV_CTRL_2_70 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_71 = zz_zz_decode_ENV_CTRL_2_72));
  zz_zz_decode_ENV_CTRL_2_75 <= pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_76) = pkg_stdLogicVector("00000000000000000000000000100000"));
  zz_zz_decode_ENV_CTRL_2_79 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_80 = zz_zz_decode_ENV_CTRL_2_81));
  zz_zz_decode_ENV_CTRL_2_82 <= pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_83),pkg_cat(zz_zz_decode_ENV_CTRL_2_85,zz_zz_decode_ENV_CTRL_2_88));
  zz_zz_decode_ENV_CTRL_2_92 <= pkg_toStdLogicVector(zz_decode_ENV_CTRL_5);
  zz_zz_decode_ENV_CTRL_2_93 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_94 = zz_zz_decode_ENV_CTRL_2_95));
  zz_zz_decode_ENV_CTRL_2_97 <= pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_5),pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_98));
  zz_zz_decode_ENV_CTRL_2_100 <= pkg_stdLogicVector("00");
  zz_zz_decode_ENV_CTRL_2_101 <= pkg_toStdLogic(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_102) /= pkg_stdLogicVector("0"));
  zz_zz_decode_ENV_CTRL_2_104 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_105 /= zz_zz_decode_ENV_CTRL_2_108));
  zz_zz_decode_ENV_CTRL_2_109 <= pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_110),pkg_cat(zz_zz_decode_ENV_CTRL_2_116,zz_zz_decode_ENV_CTRL_2_120));
  zz_zz_decode_ENV_CTRL_2_68 <= pkg_stdLogicVector("00000000000000000100000000100000");
  zz_zz_decode_ENV_CTRL_2_71 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000010000000000000000000100000"));
  zz_zz_decode_ENV_CTRL_2_72 <= pkg_stdLogicVector("00000000000000000000000000100000");
  zz_zz_decode_ENV_CTRL_2_76 <= pkg_stdLogicVector("00000010000000000000000001100000");
  zz_zz_decode_ENV_CTRL_2_80 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000001000000010000"));
  zz_zz_decode_ENV_CTRL_2_81 <= pkg_stdLogicVector("00000000000000000001000000010000");
  zz_zz_decode_ENV_CTRL_2_83 <= pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_84) = pkg_stdLogicVector("00000000000000000010000000010000"));
  zz_zz_decode_ENV_CTRL_2_85 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_86 = zz_zz_decode_ENV_CTRL_2_87));
  zz_zz_decode_ENV_CTRL_2_88 <= pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_89),pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_90));
  zz_zz_decode_ENV_CTRL_2_94 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001110000"));
  zz_zz_decode_ENV_CTRL_2_95 <= pkg_stdLogicVector("00000000000000000000000000100000");
  zz_zz_decode_ENV_CTRL_2_98 <= pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_99) = pkg_stdLogicVector("00000000000000000000000000000000"));
  zz_zz_decode_ENV_CTRL_2_102 <= pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_103) = pkg_stdLogicVector("00000000000000000100000000010000"));
  zz_zz_decode_ENV_CTRL_2_105 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_106 = zz_zz_decode_ENV_CTRL_2_107));
  zz_zz_decode_ENV_CTRL_2_108 <= pkg_stdLogicVector("0");
  zz_zz_decode_ENV_CTRL_2_110 <= pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_111,zz_zz_decode_ENV_CTRL_2_113) /= pkg_stdLogicVector("0000"));
  zz_zz_decode_ENV_CTRL_2_116 <= pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_117 /= zz_zz_decode_ENV_CTRL_2_119));
  zz_zz_decode_ENV_CTRL_2_120 <= pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_121),pkg_cat(zz_zz_decode_ENV_CTRL_2_127,zz_zz_decode_ENV_CTRL_2_131));
  zz_zz_decode_ENV_CTRL_2_84 <= pkg_stdLogicVector("00000000000000000010000000010000");
  zz_zz_decode_ENV_CTRL_2_86 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001010000"));
  zz_zz_decode_ENV_CTRL_2_87 <= pkg_stdLogicVector("00000000000000000000000000010000");
  zz_zz_decode_ENV_CTRL_2_89 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000001100")) = pkg_stdLogicVector("00000000000000000000000000000100"));
  zz_zz_decode_ENV_CTRL_2_90 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000101000")) = pkg_stdLogicVector("00000000000000000000000000000000"));
  zz_zz_decode_ENV_CTRL_2_99 <= pkg_stdLogicVector("00000000000000000000000000100000");
  zz_zz_decode_ENV_CTRL_2_103 <= pkg_stdLogicVector("00000000000000000100000000010100");
  zz_zz_decode_ENV_CTRL_2_106 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000110000000010100"));
  zz_zz_decode_ENV_CTRL_2_107 <= pkg_stdLogicVector("00000000000000000010000000010000");
  zz_zz_decode_ENV_CTRL_2_111 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_112) = pkg_stdLogicVector("00000000000000000000000000000000")));
  zz_zz_decode_ENV_CTRL_2_113 <= pkg_cat(pkg_toStdLogicVector(zz_decode_ENV_CTRL_4),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_114),pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_115)));
  zz_zz_decode_ENV_CTRL_2_117 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_118) = pkg_stdLogicVector("00000000000000000000000000000000")));
  zz_zz_decode_ENV_CTRL_2_119 <= pkg_stdLogicVector("0");
  zz_zz_decode_ENV_CTRL_2_121 <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_122),pkg_cat(zz_zz_decode_ENV_CTRL_2_123,zz_zz_decode_ENV_CTRL_2_125)) /= pkg_stdLogicVector("000"));
  zz_zz_decode_ENV_CTRL_2_127 <= pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_128,zz_zz_decode_ENV_CTRL_2_130) /= pkg_stdLogicVector("00")));
  zz_zz_decode_ENV_CTRL_2_131 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_132 /= zz_zz_decode_ENV_CTRL_2_135)),pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_136 /= zz_zz_decode_ENV_CTRL_2_138)));
  zz_zz_decode_ENV_CTRL_2_112 <= pkg_stdLogicVector("00000000000000000000000001000100");
  zz_zz_decode_ENV_CTRL_2_114 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000110000000000100")) = pkg_stdLogicVector("00000000000000000010000000000000"));
  zz_zz_decode_ENV_CTRL_2_115 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000101000000000100")) = pkg_stdLogicVector("00000000000000000001000000000000"));
  zz_zz_decode_ENV_CTRL_2_118 <= pkg_stdLogicVector("00000000000000000000000001011000");
  zz_zz_decode_ENV_CTRL_2_122 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001000100")) = pkg_stdLogicVector("00000000000000000000000001000000"));
  zz_zz_decode_ENV_CTRL_2_123 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_124) = pkg_stdLogicVector("00000000000000000010000000010000")));
  zz_zz_decode_ENV_CTRL_2_125 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_126) = pkg_stdLogicVector("01000000000000000000000000110000")));
  zz_zz_decode_ENV_CTRL_2_128 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_129) = pkg_stdLogicVector("00000000000000000000000000000100")));
  zz_zz_decode_ENV_CTRL_2_130 <= pkg_toStdLogicVector(zz_decode_ENV_CTRL_3);
  zz_zz_decode_ENV_CTRL_2_132 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_133 = zz_zz_decode_ENV_CTRL_2_134)),pkg_toStdLogicVector(zz_decode_ENV_CTRL_3));
  zz_zz_decode_ENV_CTRL_2_135 <= pkg_stdLogicVector("00");
  zz_zz_decode_ENV_CTRL_2_136 <= pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2_137) = pkg_stdLogicVector("00000000000000000001000000001000")));
  zz_zz_decode_ENV_CTRL_2_138 <= pkg_stdLogicVector("0");
  zz_zz_decode_ENV_CTRL_2_124 <= pkg_stdLogicVector("00000000000000000010000000010100");
  zz_zz_decode_ENV_CTRL_2_126 <= pkg_stdLogicVector("01000000000000000000000000110100");
  zz_zz_decode_ENV_CTRL_2_129 <= pkg_stdLogicVector("00000000000000000000000000010100");
  zz_zz_decode_ENV_CTRL_2_133 <= (decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001000100"));
  zz_zz_decode_ENV_CTRL_2_134 <= pkg_stdLogicVector("00000000000000000000000000000100");
  zz_zz_decode_ENV_CTRL_2_137 <= pkg_stdLogicVector("00000000000000000101000001001000");
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_2 = '1' then
        IBusCachedPlugin_predictor_history(to_integer(IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_address)) <= zz_IBusCachedPlugin_predictor_history_port;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if IBusCachedPlugin_iBusRsp_stages_0_output_ready = '1' then
        zz_IBusCachedPlugin_predictor_history_port0 <= IBusCachedPlugin_predictor_history(to_integer(zz_zz_IBusCachedPlugin_predictor_buffer_line_source_1));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_decode_RegFilePlugin_rs1Data = '1' then
        zz_RegFilePlugin_regFile_port0 <= RegFilePlugin_regFile(to_integer(decode_RegFilePlugin_regFileReadAddress1));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_decode_RegFilePlugin_rs2Data = '1' then
        zz_RegFilePlugin_regFile_port0_1 <= RegFilePlugin_regFile(to_integer(decode_RegFilePlugin_regFileReadAddress2));
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if zz_1 = '1' then
        RegFilePlugin_regFile(to_integer(lastStageRegFileWrite_payload_address)) <= lastStageRegFileWrite_payload_data;
      end if;
    end if;
  end process;

  IBusCachedPlugin_cache : entity work.InstructionCache
    port map ( 
      io_flush => IBusCachedPlugin_cache_io_flush,
      io_cpu_prefetch_isValid => IBusCachedPlugin_cache_io_cpu_prefetch_isValid,
      io_cpu_prefetch_haltIt => IBusCachedPlugin_cache_io_cpu_prefetch_haltIt,
      io_cpu_prefetch_pc => IBusCachedPlugin_iBusRsp_stages_0_input_payload,
      io_cpu_fetch_isValid => IBusCachedPlugin_cache_io_cpu_fetch_isValid,
      io_cpu_fetch_isStuck => IBusCachedPlugin_cache_io_cpu_fetch_isStuck,
      io_cpu_fetch_isRemoved => IBusCachedPlugin_cache_io_cpu_fetch_isRemoved,
      io_cpu_fetch_pc => IBusCachedPlugin_iBusRsp_stages_1_input_payload,
      io_cpu_fetch_data => IBusCachedPlugin_cache_io_cpu_fetch_data,
      io_cpu_fetch_mmuRsp_physicalAddress => IBusCachedPlugin_mmuBus_rsp_physicalAddress,
      io_cpu_fetch_mmuRsp_isIoAccess => IBusCachedPlugin_mmuBus_rsp_isIoAccess,
      io_cpu_fetch_mmuRsp_isPaging => IBusCachedPlugin_mmuBus_rsp_isPaging,
      io_cpu_fetch_mmuRsp_allowRead => IBusCachedPlugin_mmuBus_rsp_allowRead,
      io_cpu_fetch_mmuRsp_allowWrite => IBusCachedPlugin_mmuBus_rsp_allowWrite,
      io_cpu_fetch_mmuRsp_allowExecute => IBusCachedPlugin_mmuBus_rsp_allowExecute,
      io_cpu_fetch_mmuRsp_exception => IBusCachedPlugin_mmuBus_rsp_exception,
      io_cpu_fetch_mmuRsp_refilling => IBusCachedPlugin_mmuBus_rsp_refilling,
      io_cpu_fetch_mmuRsp_bypassTranslation => IBusCachedPlugin_mmuBus_rsp_bypassTranslation,
      io_cpu_fetch_physicalAddress => IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress,
      io_cpu_decode_isValid => IBusCachedPlugin_cache_io_cpu_decode_isValid,
      io_cpu_decode_isStuck => IBusCachedPlugin_cache_io_cpu_decode_isStuck,
      io_cpu_decode_pc => IBusCachedPlugin_iBusRsp_stages_2_input_payload,
      io_cpu_decode_physicalAddress => IBusCachedPlugin_cache_io_cpu_decode_physicalAddress,
      io_cpu_decode_data => IBusCachedPlugin_cache_io_cpu_decode_data,
      io_cpu_decode_cacheMiss => IBusCachedPlugin_cache_io_cpu_decode_cacheMiss,
      io_cpu_decode_error => IBusCachedPlugin_cache_io_cpu_decode_error,
      io_cpu_decode_mmuRefilling => IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling,
      io_cpu_decode_mmuException => IBusCachedPlugin_cache_io_cpu_decode_mmuException,
      io_cpu_decode_isUser => IBusCachedPlugin_cache_io_cpu_decode_isUser,
      io_cpu_fill_valid => IBusCachedPlugin_cache_io_cpu_fill_valid,
      io_cpu_fill_payload => IBusCachedPlugin_cache_io_cpu_decode_physicalAddress,
      io_mem_cmd_valid => IBusCachedPlugin_cache_io_mem_cmd_valid,
      io_mem_cmd_ready => iBus_cmd_ready,
      io_mem_cmd_payload_address => IBusCachedPlugin_cache_io_mem_cmd_payload_address,
      io_mem_cmd_payload_size => IBusCachedPlugin_cache_io_mem_cmd_payload_size,
      io_mem_rsp_valid => iBus_rsp_valid,
      io_mem_rsp_payload_data => iBus_rsp_payload_data,
      io_mem_rsp_payload_error => iBus_rsp_payload_error,
      zz_when_Fetcher_l398 => switch_Fetcher_l362,
      zz_io_cpu_fetch_data_regNextWhen => IBusCachedPlugin_injectionPort_payload,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  dataCache_1 : entity work.DataCache
    port map ( 
      io_cpu_execute_isValid => dataCache_1_io_cpu_execute_isValid,
      io_cpu_execute_address => dataCache_1_io_cpu_execute_address,
      io_cpu_execute_haltIt => dataCache_1_io_cpu_execute_haltIt,
      io_cpu_execute_args_wr => execute_MEMORY_WR,
      io_cpu_execute_args_size => execute_DBusCachedPlugin_size,
      io_cpu_execute_args_totalyConsistent => execute_MEMORY_FORCE_CONSTISTENCY,
      io_cpu_execute_refilling => dataCache_1_io_cpu_execute_refilling,
      io_cpu_memory_isValid => dataCache_1_io_cpu_memory_isValid,
      io_cpu_memory_isStuck => memory_arbitration_isStuck,
      io_cpu_memory_isWrite => dataCache_1_io_cpu_memory_isWrite,
      io_cpu_memory_address => dataCache_1_io_cpu_memory_address,
      io_cpu_memory_mmuRsp_physicalAddress => DBusCachedPlugin_mmuBus_rsp_physicalAddress,
      io_cpu_memory_mmuRsp_isIoAccess => dataCache_1_io_cpu_memory_mmuRsp_isIoAccess,
      io_cpu_memory_mmuRsp_isPaging => DBusCachedPlugin_mmuBus_rsp_isPaging,
      io_cpu_memory_mmuRsp_allowRead => DBusCachedPlugin_mmuBus_rsp_allowRead,
      io_cpu_memory_mmuRsp_allowWrite => DBusCachedPlugin_mmuBus_rsp_allowWrite,
      io_cpu_memory_mmuRsp_allowExecute => DBusCachedPlugin_mmuBus_rsp_allowExecute,
      io_cpu_memory_mmuRsp_exception => DBusCachedPlugin_mmuBus_rsp_exception,
      io_cpu_memory_mmuRsp_refilling => DBusCachedPlugin_mmuBus_rsp_refilling,
      io_cpu_memory_mmuRsp_bypassTranslation => DBusCachedPlugin_mmuBus_rsp_bypassTranslation,
      io_cpu_writeBack_isValid => dataCache_1_io_cpu_writeBack_isValid,
      io_cpu_writeBack_isStuck => writeBack_arbitration_isStuck,
      io_cpu_writeBack_isUser => dataCache_1_io_cpu_writeBack_isUser,
      io_cpu_writeBack_haltIt => dataCache_1_io_cpu_writeBack_haltIt,
      io_cpu_writeBack_isWrite => dataCache_1_io_cpu_writeBack_isWrite,
      io_cpu_writeBack_storeData => dataCache_1_io_cpu_writeBack_storeData,
      io_cpu_writeBack_data => dataCache_1_io_cpu_writeBack_data,
      io_cpu_writeBack_address => dataCache_1_io_cpu_writeBack_address,
      io_cpu_writeBack_mmuException => dataCache_1_io_cpu_writeBack_mmuException,
      io_cpu_writeBack_unalignedAccess => dataCache_1_io_cpu_writeBack_unalignedAccess,
      io_cpu_writeBack_accessError => dataCache_1_io_cpu_writeBack_accessError,
      io_cpu_writeBack_keepMemRspData => dataCache_1_io_cpu_writeBack_keepMemRspData,
      io_cpu_writeBack_fence_SW => dataCache_1_io_cpu_writeBack_fence_SW,
      io_cpu_writeBack_fence_SR => dataCache_1_io_cpu_writeBack_fence_SR,
      io_cpu_writeBack_fence_SO => dataCache_1_io_cpu_writeBack_fence_SO,
      io_cpu_writeBack_fence_SI => dataCache_1_io_cpu_writeBack_fence_SI,
      io_cpu_writeBack_fence_PW => dataCache_1_io_cpu_writeBack_fence_PW,
      io_cpu_writeBack_fence_PR => dataCache_1_io_cpu_writeBack_fence_PR,
      io_cpu_writeBack_fence_PO => dataCache_1_io_cpu_writeBack_fence_PO,
      io_cpu_writeBack_fence_PI => dataCache_1_io_cpu_writeBack_fence_PI,
      io_cpu_writeBack_fence_FM => dataCache_1_io_cpu_writeBack_fence_FM,
      io_cpu_writeBack_exclusiveOk => dataCache_1_io_cpu_writeBack_exclusiveOk,
      io_cpu_redo => dataCache_1_io_cpu_redo,
      io_cpu_flush_valid => dataCache_1_io_cpu_flush_valid,
      io_cpu_flush_ready => dataCache_1_io_cpu_flush_ready,
      io_mem_cmd_valid => dataCache_1_io_mem_cmd_valid,
      io_mem_cmd_ready => dBus_cmd_ready,
      io_mem_cmd_payload_wr => dataCache_1_io_mem_cmd_payload_wr,
      io_mem_cmd_payload_uncached => dataCache_1_io_mem_cmd_payload_uncached,
      io_mem_cmd_payload_address => dataCache_1_io_mem_cmd_payload_address,
      io_mem_cmd_payload_data => dataCache_1_io_mem_cmd_payload_data,
      io_mem_cmd_payload_mask => dataCache_1_io_mem_cmd_payload_mask,
      io_mem_cmd_payload_size => dataCache_1_io_mem_cmd_payload_size,
      io_mem_cmd_payload_last => dataCache_1_io_mem_cmd_payload_last,
      io_mem_rsp_valid => dBus_rsp_valid,
      io_mem_rsp_payload_last => dBus_rsp_payload_last,
      io_mem_rsp_payload_data => dBus_rsp_payload_data,
      io_mem_rsp_payload_error => dBus_rsp_payload_error,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  process(zz_IBusCachedPlugin_jump_pcLoad_payload_5,DBusCachedPlugin_redoBranch_payload,CsrPlugin_jumpInterface_payload,BranchPlugin_jumpInterface_payload)
  begin
    case zz_IBusCachedPlugin_jump_pcLoad_payload_5 is
      when "00" =>
        zz_IBusCachedPlugin_jump_pcLoad_payload_4 <= DBusCachedPlugin_redoBranch_payload;
      when "01" =>
        zz_IBusCachedPlugin_jump_pcLoad_payload_4 <= CsrPlugin_jumpInterface_payload;
      when others =>
        zz_IBusCachedPlugin_jump_pcLoad_payload_4 <= BranchPlugin_jumpInterface_payload;
    end case;
  end process;

  process(zz_writeBack_DBusCachedPlugin_rspShifted_1,writeBack_DBusCachedPlugin_rspSplits_0,writeBack_DBusCachedPlugin_rspSplits_1,writeBack_DBusCachedPlugin_rspSplits_2,writeBack_DBusCachedPlugin_rspSplits_3)
  begin
    case zz_writeBack_DBusCachedPlugin_rspShifted_1 is
      when "00" =>
        zz_writeBack_DBusCachedPlugin_rspShifted <= writeBack_DBusCachedPlugin_rspSplits_0;
      when "01" =>
        zz_writeBack_DBusCachedPlugin_rspShifted <= writeBack_DBusCachedPlugin_rspSplits_1;
      when "10" =>
        zz_writeBack_DBusCachedPlugin_rspShifted <= writeBack_DBusCachedPlugin_rspSplits_2;
      when others =>
        zz_writeBack_DBusCachedPlugin_rspShifted <= writeBack_DBusCachedPlugin_rspSplits_3;
    end case;
  end process;

  process(zz_writeBack_DBusCachedPlugin_rspShifted_3,writeBack_DBusCachedPlugin_rspSplits_1,writeBack_DBusCachedPlugin_rspSplits_3)
  begin
    case zz_writeBack_DBusCachedPlugin_rspShifted_3 is
      when "0" =>
        zz_writeBack_DBusCachedPlugin_rspShifted_2 <= writeBack_DBusCachedPlugin_rspSplits_1;
      when others =>
        zz_writeBack_DBusCachedPlugin_rspShifted_2 <= writeBack_DBusCachedPlugin_rspSplits_3;
    end case;
  end process;

  memory_MUL_LOW <= (((pkg_signed("0000000000000000000000000000000000000000000000000000") + pkg_resize(signed(pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(false)),std_logic_vector(memory_MUL_LL))),52)) + pkg_resize(pkg_shiftLeft(memory_MUL_LH,16),52)) + pkg_resize(pkg_shiftLeft(memory_MUL_HL,16),52));
  execute_TARGET_MISSMATCH2 <= pkg_toStdLogic(decode_PC /= execute_BRANCH_CALC);
  execute_NEXT_PC2 <= (execute_PC + pkg_unsigned("00000000000000000000000000000100"));
  execute_BRANCH_DO <= zz_execute_BRANCH_DO_1;
  memory_MUL_HH <= execute_to_memory_MUL_HH;
  execute_MUL_HH <= (execute_MulPlugin_aHigh * execute_MulPlugin_bHigh);
  execute_MUL_HL <= (execute_MulPlugin_aHigh * execute_MulPlugin_bSLow);
  execute_MUL_LH <= (execute_MulPlugin_aSLow * execute_MulPlugin_bHigh);
  execute_MUL_LL <= (execute_MulPlugin_aULow * execute_MulPlugin_bULow);
  execute_REGFILE_WRITE_DATA <= zz_execute_REGFILE_WRITE_DATA;
  memory_MEMORY_STORE_DATA_RF <= execute_to_memory_MEMORY_STORE_DATA_RF;
  execute_MEMORY_STORE_DATA_RF <= zz_execute_MEMORY_STORE_DATA_RF;
  decode_DO_EBREAK <= (((not DebugPlugin_haltIt) and (decode_IS_EBREAK or pkg_toStdLogic(false))) and DebugPlugin_allowEBreak);
  decode_CSR_READ_OPCODE <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,13,7) /= pkg_stdLogicVector("0100000"));
  decode_CSR_WRITE_OPCODE <= (not ((pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,14,13) = pkg_stdLogicVector("01")) and pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,19,15) = pkg_stdLogicVector("00000"))) or (pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,14,13) = pkg_stdLogicVector("11")) and pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,19,15) = pkg_stdLogicVector("00000")))));
  decode_SRC2_FORCE_ZERO <= (decode_SRC_ADD_ZERO and (not decode_SRC_USE_SUB_LESS));
  zz_memory_to_writeBack_ENV_CTRL <= zz_memory_to_writeBack_ENV_CTRL_1;
  zz_execute_to_memory_ENV_CTRL <= zz_execute_to_memory_ENV_CTRL_1;
  decode_ENV_CTRL <= zz_decode_ENV_CTRL;
  zz_decode_to_execute_ENV_CTRL <= zz_decode_to_execute_ENV_CTRL_1;
  decode_IS_CSR <= pkg_extract(zz_decode_ENV_CTRL_2,29);
  decode_BRANCH_CTRL <= zz_decode_BRANCH_CTRL;
  zz_decode_to_execute_BRANCH_CTRL <= zz_decode_to_execute_BRANCH_CTRL_1;
  decode_IS_RS2_SIGNED <= pkg_extract(zz_decode_ENV_CTRL_2,26);
  decode_IS_RS1_SIGNED <= pkg_extract(zz_decode_ENV_CTRL_2,25);
  decode_IS_DIV <= pkg_extract(zz_decode_ENV_CTRL_2,24);
  memory_IS_MUL <= execute_to_memory_IS_MUL;
  execute_IS_MUL <= decode_to_execute_IS_MUL;
  decode_IS_MUL <= pkg_extract(zz_decode_ENV_CTRL_2,23);
  decode_SHIFT_CTRL <= zz_decode_SHIFT_CTRL;
  zz_decode_to_execute_SHIFT_CTRL <= zz_decode_to_execute_SHIFT_CTRL_1;
  decode_ALU_BITWISE_CTRL <= zz_decode_ALU_BITWISE_CTRL;
  zz_decode_to_execute_ALU_BITWISE_CTRL <= zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  decode_SRC_LESS_UNSIGNED <= pkg_extract(zz_decode_ENV_CTRL_2,17);
  decode_MEMORY_MANAGMENT <= pkg_extract(zz_decode_ENV_CTRL_2,16);
  memory_MEMORY_WR <= execute_to_memory_MEMORY_WR;
  decode_MEMORY_WR <= pkg_extract(zz_decode_ENV_CTRL_2,13);
  execute_BYPASSABLE_MEMORY_STAGE <= decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  decode_BYPASSABLE_MEMORY_STAGE <= pkg_extract(zz_decode_ENV_CTRL_2,12);
  decode_BYPASSABLE_EXECUTE_STAGE <= pkg_extract(zz_decode_ENV_CTRL_2,11);
  decode_SRC2_CTRL <= zz_decode_SRC2_CTRL;
  zz_decode_to_execute_SRC2_CTRL <= zz_decode_to_execute_SRC2_CTRL_1;
  decode_ALU_CTRL <= zz_decode_ALU_CTRL;
  zz_decode_to_execute_ALU_CTRL <= zz_decode_to_execute_ALU_CTRL_1;
  decode_SRC1_CTRL <= zz_decode_SRC1_CTRL;
  zz_decode_to_execute_SRC1_CTRL <= zz_decode_to_execute_SRC1_CTRL_1;
  decode_MEMORY_FORCE_CONSTISTENCY <= pkg_toStdLogic(false);
  execute_PREDICTION_CONTEXT_hazard <= decode_to_execute_PREDICTION_CONTEXT_hazard;
  execute_PREDICTION_CONTEXT_hit <= decode_to_execute_PREDICTION_CONTEXT_hit;
  execute_PREDICTION_CONTEXT_line_source <= decode_to_execute_PREDICTION_CONTEXT_line_source;
  execute_PREDICTION_CONTEXT_line_branchWish <= decode_to_execute_PREDICTION_CONTEXT_line_branchWish;
  execute_PREDICTION_CONTEXT_line_target <= decode_to_execute_PREDICTION_CONTEXT_line_target;
  decode_PREDICTION_CONTEXT_hazard <= IBusCachedPlugin_predictor_injectorContext_hazard;
  decode_PREDICTION_CONTEXT_hit <= IBusCachedPlugin_predictor_injectorContext_hit;
  decode_PREDICTION_CONTEXT_line_source <= IBusCachedPlugin_predictor_injectorContext_line_source;
  decode_PREDICTION_CONTEXT_line_branchWish <= IBusCachedPlugin_predictor_injectorContext_line_branchWish;
  decode_PREDICTION_CONTEXT_line_target <= IBusCachedPlugin_predictor_injectorContext_line_target;
  writeBack_FORMAL_PC_NEXT <= memory_to_writeBack_FORMAL_PC_NEXT;
  memory_FORMAL_PC_NEXT <= execute_to_memory_FORMAL_PC_NEXT;
  execute_FORMAL_PC_NEXT <= decode_to_execute_FORMAL_PC_NEXT;
  decode_FORMAL_PC_NEXT <= (decode_PC + pkg_unsigned("00000000000000000000000000000100"));
  execute_DO_EBREAK <= decode_to_execute_DO_EBREAK;
  decode_IS_EBREAK <= pkg_extract(zz_decode_ENV_CTRL_2,31);
  execute_CSR_READ_OPCODE <= decode_to_execute_CSR_READ_OPCODE;
  execute_CSR_WRITE_OPCODE <= decode_to_execute_CSR_WRITE_OPCODE;
  execute_IS_CSR <= decode_to_execute_IS_CSR;
  memory_ENV_CTRL <= zz_memory_ENV_CTRL;
  execute_ENV_CTRL <= zz_execute_ENV_CTRL;
  writeBack_ENV_CTRL <= zz_writeBack_ENV_CTRL;
  memory_NEXT_PC2 <= execute_to_memory_NEXT_PC2;
  memory_PC <= execute_to_memory_PC;
  memory_BRANCH_CALC <= execute_to_memory_BRANCH_CALC;
  memory_TARGET_MISSMATCH2 <= execute_to_memory_TARGET_MISSMATCH2;
  memory_BRANCH_DO <= execute_to_memory_BRANCH_DO;
  execute_BRANCH_CALC <= unsigned(pkg_cat(std_logic_vector(pkg_extract(execute_BranchPlugin_branchAdder,31,1)),std_logic_vector(pkg_unsigned("0"))));
  execute_BRANCH_SRC22 <= unsigned(zz_execute_BRANCH_SRC22_6);
  execute_PC <= decode_to_execute_PC;
  execute_BRANCH_CTRL <= zz_execute_BRANCH_CTRL;
  decode_RS2_USE <= pkg_extract(zz_decode_ENV_CTRL_2,15);
  decode_RS1_USE <= pkg_extract(zz_decode_ENV_CTRL_2,5);
  execute_REGFILE_WRITE_VALID <= decode_to_execute_REGFILE_WRITE_VALID;
  execute_BYPASSABLE_EXECUTE_STAGE <= decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  memory_REGFILE_WRITE_VALID <= execute_to_memory_REGFILE_WRITE_VALID;
  memory_BYPASSABLE_MEMORY_STAGE <= execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  writeBack_REGFILE_WRITE_VALID <= memory_to_writeBack_REGFILE_WRITE_VALID;
  process(decode_RegFilePlugin_rs2Data,HazardSimplePlugin_writeBackBuffer_valid,HazardSimplePlugin_addr1Match,HazardSimplePlugin_writeBackBuffer_payload_data,when_HazardSimplePlugin_l45,when_HazardSimplePlugin_l47,when_HazardSimplePlugin_l51,zz_decode_RS2_2,when_HazardSimplePlugin_l45_1,memory_BYPASSABLE_MEMORY_STAGE,when_HazardSimplePlugin_l51_1,zz_decode_RS2,when_HazardSimplePlugin_l45_2,execute_BYPASSABLE_EXECUTE_STAGE,when_HazardSimplePlugin_l51_2,zz_decode_RS2_1)
  begin
    decode_RS2 <= decode_RegFilePlugin_rs2Data;
    if HazardSimplePlugin_writeBackBuffer_valid = '1' then
      if HazardSimplePlugin_addr1Match = '1' then
        decode_RS2 <= HazardSimplePlugin_writeBackBuffer_payload_data;
      end if;
    end if;
    if when_HazardSimplePlugin_l45 = '1' then
      if when_HazardSimplePlugin_l47 = '1' then
        if when_HazardSimplePlugin_l51 = '1' then
          decode_RS2 <= zz_decode_RS2_2;
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l45_1 = '1' then
      if memory_BYPASSABLE_MEMORY_STAGE = '1' then
        if when_HazardSimplePlugin_l51_1 = '1' then
          decode_RS2 <= zz_decode_RS2;
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l45_2 = '1' then
      if execute_BYPASSABLE_EXECUTE_STAGE = '1' then
        if when_HazardSimplePlugin_l51_2 = '1' then
          decode_RS2 <= zz_decode_RS2_1;
        end if;
      end if;
    end if;
  end process;

  process(decode_RegFilePlugin_rs1Data,HazardSimplePlugin_writeBackBuffer_valid,HazardSimplePlugin_addr0Match,HazardSimplePlugin_writeBackBuffer_payload_data,when_HazardSimplePlugin_l45,when_HazardSimplePlugin_l47,when_HazardSimplePlugin_l48,zz_decode_RS2_2,when_HazardSimplePlugin_l45_1,memory_BYPASSABLE_MEMORY_STAGE,when_HazardSimplePlugin_l48_1,zz_decode_RS2,when_HazardSimplePlugin_l45_2,execute_BYPASSABLE_EXECUTE_STAGE,when_HazardSimplePlugin_l48_2,zz_decode_RS2_1)
  begin
    decode_RS1 <= decode_RegFilePlugin_rs1Data;
    if HazardSimplePlugin_writeBackBuffer_valid = '1' then
      if HazardSimplePlugin_addr0Match = '1' then
        decode_RS1 <= HazardSimplePlugin_writeBackBuffer_payload_data;
      end if;
    end if;
    if when_HazardSimplePlugin_l45 = '1' then
      if when_HazardSimplePlugin_l47 = '1' then
        if when_HazardSimplePlugin_l48 = '1' then
          decode_RS1 <= zz_decode_RS2_2;
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l45_1 = '1' then
      if memory_BYPASSABLE_MEMORY_STAGE = '1' then
        if when_HazardSimplePlugin_l48_1 = '1' then
          decode_RS1 <= zz_decode_RS2;
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l45_2 = '1' then
      if execute_BYPASSABLE_EXECUTE_STAGE = '1' then
        if when_HazardSimplePlugin_l48_2 = '1' then
          decode_RS1 <= zz_decode_RS2_1;
        end if;
      end if;
    end if;
  end process;

  execute_IS_RS1_SIGNED <= decode_to_execute_IS_RS1_SIGNED;
  execute_IS_DIV <= decode_to_execute_IS_DIV;
  execute_IS_RS2_SIGNED <= decode_to_execute_IS_RS2_SIGNED;
  process(memory_REGFILE_WRITE_DATA,when_MulDivIterativePlugin_l128,memory_DivPlugin_div_result)
  begin
    zz_decode_RS2 <= memory_REGFILE_WRITE_DATA;
    if when_MulDivIterativePlugin_l128 = '1' then
      zz_decode_RS2 <= memory_DivPlugin_div_result;
    end if;
  end process;

  memory_INSTRUCTION <= execute_to_memory_INSTRUCTION;
  memory_IS_DIV <= execute_to_memory_IS_DIV;
  writeBack_IS_MUL <= memory_to_writeBack_IS_MUL;
  writeBack_MUL_HH <= memory_to_writeBack_MUL_HH;
  writeBack_MUL_LOW <= memory_to_writeBack_MUL_LOW;
  memory_MUL_HL <= execute_to_memory_MUL_HL;
  memory_MUL_LH <= execute_to_memory_MUL_LH;
  memory_MUL_LL <= execute_to_memory_MUL_LL;
  execute_RS1 <= decode_to_execute_RS1;
  execute_SHIFT_RIGHT <= std_logic_vector(pkg_extract(pkg_shiftRight(signed(pkg_cat(pkg_toStdLogicVector((pkg_toStdLogic(execute_SHIFT_CTRL = ShiftCtrlEnum_seq_SRA_1) and pkg_extract(execute_FullBarrelShifterPlugin_reversed,31))),execute_FullBarrelShifterPlugin_reversed)),execute_FullBarrelShifterPlugin_amplitude),31,0));
  process(execute_REGFILE_WRITE_DATA,execute_arbitration_isValid,execute_SHIFT_CTRL,zz_decode_RS2_3,execute_SHIFT_RIGHT,when_CsrPlugin_l1176,CsrPlugin_csrMapping_readDataSignal)
  begin
    zz_decode_RS2_1 <= execute_REGFILE_WRITE_DATA;
    if execute_arbitration_isValid = '1' then
      case execute_SHIFT_CTRL is
        when ShiftCtrlEnum_seq_SLL_1 =>
          zz_decode_RS2_1 <= zz_decode_RS2_3;
        when ShiftCtrlEnum_seq_SRL_1 | ShiftCtrlEnum_seq_SRA_1 =>
          zz_decode_RS2_1 <= execute_SHIFT_RIGHT;
        when others =>
      end case;
    end if;
    if when_CsrPlugin_l1176 = '1' then
      zz_decode_RS2_1 <= CsrPlugin_csrMapping_readDataSignal;
    end if;
  end process;

  execute_SHIFT_CTRL <= zz_execute_SHIFT_CTRL;
  execute_SRC_LESS_UNSIGNED <= decode_to_execute_SRC_LESS_UNSIGNED;
  execute_SRC2_FORCE_ZERO <= decode_to_execute_SRC2_FORCE_ZERO;
  execute_SRC_USE_SUB_LESS <= decode_to_execute_SRC_USE_SUB_LESS;
  zz_execute_SRC2 <= execute_PC;
  execute_SRC2_CTRL <= zz_execute_SRC2_CTRL;
  execute_SRC1_CTRL <= zz_execute_SRC1_CTRL;
  decode_SRC_USE_SUB_LESS <= pkg_extract(zz_decode_ENV_CTRL_2,3);
  decode_SRC_ADD_ZERO <= pkg_extract(zz_decode_ENV_CTRL_2,20);
  execute_SRC_ADD_SUB <= execute_SrcPlugin_addSub;
  execute_SRC_LESS <= execute_SrcPlugin_less;
  execute_ALU_CTRL <= zz_execute_ALU_CTRL;
  execute_SRC2 <= zz_execute_SRC2_5;
  execute_SRC1 <= zz_execute_SRC1;
  execute_ALU_BITWISE_CTRL <= zz_execute_ALU_BITWISE_CTRL;
  zz_lastStageRegFileWrite_payload_address <= writeBack_INSTRUCTION;
  zz_lastStageRegFileWrite_valid <= writeBack_REGFILE_WRITE_VALID;
  process(lastStageRegFileWrite_valid)
  begin
    zz_1 <= pkg_toStdLogic(false);
    if lastStageRegFileWrite_valid = '1' then
      zz_1 <= pkg_toStdLogic(true);
    end if;
  end process;

  decode_INSTRUCTION_ANTICIPATED <= pkg_mux(decode_arbitration_isStuck,decode_INSTRUCTION,IBusCachedPlugin_cache_io_cpu_fetch_data);
  process(zz_decode_ENV_CTRL_2,when_RegFilePlugin_l63)
  begin
    decode_REGFILE_WRITE_VALID <= pkg_extract(zz_decode_ENV_CTRL_2,10);
    if when_RegFilePlugin_l63 = '1' then
      decode_REGFILE_WRITE_VALID <= pkg_toStdLogic(false);
    end if;
  end process;

  decode_LEGAL_INSTRUCTION <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001011111")) = pkg_stdLogicVector("00000000000000000000000000010111"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001111111")) = pkg_stdLogicVector("00000000000000000000000001101111"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_decode_LEGAL_INSTRUCTION) = pkg_stdLogicVector("00000000000000000000000000000011"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_decode_LEGAL_INSTRUCTION_1 = zz_decode_LEGAL_INSTRUCTION_2)),pkg_cat(pkg_toStdLogicVector(zz_decode_LEGAL_INSTRUCTION_3),pkg_cat(zz_decode_LEGAL_INSTRUCTION_4,zz_decode_LEGAL_INSTRUCTION_5)))))) /= pkg_stdLogicVector("00000000000000000000"));
  process(writeBack_REGFILE_WRITE_DATA,when_DBusCachedPlugin_l488,writeBack_DBusCachedPlugin_rspFormated,when_MulPlugin_l147,switch_MulPlugin_l148,writeBack_MUL_LOW,writeBack_MulPlugin_result)
  begin
    zz_decode_RS2_2 <= writeBack_REGFILE_WRITE_DATA;
    if when_DBusCachedPlugin_l488 = '1' then
      zz_decode_RS2_2 <= writeBack_DBusCachedPlugin_rspFormated;
    end if;
    if when_MulPlugin_l147 = '1' then
      case switch_MulPlugin_l148 is
        when "00" =>
          zz_decode_RS2_2 <= std_logic_vector(pkg_extract(writeBack_MUL_LOW,31,0));
        when others =>
          zz_decode_RS2_2 <= std_logic_vector(pkg_extract(writeBack_MulPlugin_result,63,32));
      end case;
    end if;
  end process;

  writeBack_MEMORY_WR <= memory_to_writeBack_MEMORY_WR;
  writeBack_MEMORY_STORE_DATA_RF <= memory_to_writeBack_MEMORY_STORE_DATA_RF;
  writeBack_REGFILE_WRITE_DATA <= memory_to_writeBack_REGFILE_WRITE_DATA;
  writeBack_MEMORY_ENABLE <= memory_to_writeBack_MEMORY_ENABLE;
  memory_REGFILE_WRITE_DATA <= execute_to_memory_REGFILE_WRITE_DATA;
  memory_MEMORY_ENABLE <= execute_to_memory_MEMORY_ENABLE;
  execute_MEMORY_FORCE_CONSTISTENCY <= decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  execute_MEMORY_MANAGMENT <= decode_to_execute_MEMORY_MANAGMENT;
  execute_RS2 <= decode_to_execute_RS2;
  execute_MEMORY_WR <= decode_to_execute_MEMORY_WR;
  execute_SRC_ADD <= execute_SrcPlugin_addSub;
  execute_MEMORY_ENABLE <= decode_to_execute_MEMORY_ENABLE;
  execute_INSTRUCTION <= decode_to_execute_INSTRUCTION;
  decode_MEMORY_ENABLE <= pkg_extract(zz_decode_ENV_CTRL_2,4);
  decode_FLUSH_ALL <= pkg_extract(zz_decode_ENV_CTRL_2,0);
  process(IBusCachedPlugin_rsp_issueDetected_3,when_IBusCachedPlugin_l256)
  begin
    IBusCachedPlugin_rsp_issueDetected_4 <= IBusCachedPlugin_rsp_issueDetected_3;
    if when_IBusCachedPlugin_l256 = '1' then
      IBusCachedPlugin_rsp_issueDetected_4 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(IBusCachedPlugin_rsp_issueDetected_2,when_IBusCachedPlugin_l250)
  begin
    IBusCachedPlugin_rsp_issueDetected_3 <= IBusCachedPlugin_rsp_issueDetected_2;
    if when_IBusCachedPlugin_l250 = '1' then
      IBusCachedPlugin_rsp_issueDetected_3 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(IBusCachedPlugin_rsp_issueDetected_1,when_IBusCachedPlugin_l244)
  begin
    IBusCachedPlugin_rsp_issueDetected_2 <= IBusCachedPlugin_rsp_issueDetected_1;
    if when_IBusCachedPlugin_l244 = '1' then
      IBusCachedPlugin_rsp_issueDetected_2 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(IBusCachedPlugin_rsp_issueDetected,when_IBusCachedPlugin_l239)
  begin
    IBusCachedPlugin_rsp_issueDetected_1 <= IBusCachedPlugin_rsp_issueDetected;
    if when_IBusCachedPlugin_l239 = '1' then
      IBusCachedPlugin_rsp_issueDetected_1 <= pkg_toStdLogic(true);
    end if;
  end process;

  decode_INSTRUCTION <= IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  memory_PREDICTION_CONTEXT_hazard <= execute_to_memory_PREDICTION_CONTEXT_hazard;
  memory_PREDICTION_CONTEXT_hit <= execute_to_memory_PREDICTION_CONTEXT_hit;
  memory_PREDICTION_CONTEXT_line_source <= execute_to_memory_PREDICTION_CONTEXT_line_source;
  memory_PREDICTION_CONTEXT_line_branchWish <= execute_to_memory_PREDICTION_CONTEXT_line_branchWish;
  memory_PREDICTION_CONTEXT_line_target <= execute_to_memory_PREDICTION_CONTEXT_line_target;
  process(IBusCachedPlugin_predictor_historyWriteDelayPatched_valid)
  begin
    zz_2 <= pkg_toStdLogic(false);
    if IBusCachedPlugin_predictor_historyWriteDelayPatched_valid = '1' then
      zz_2 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(memory_FORMAL_PC_NEXT,BranchPlugin_jumpInterface_valid,BranchPlugin_jumpInterface_payload)
  begin
    zz_memory_to_writeBack_FORMAL_PC_NEXT <= memory_FORMAL_PC_NEXT;
    if BranchPlugin_jumpInterface_valid = '1' then
      zz_memory_to_writeBack_FORMAL_PC_NEXT <= BranchPlugin_jumpInterface_payload;
    end if;
  end process;

  decode_PC <= IBusCachedPlugin_iBusRsp_output_payload_pc;
  writeBack_PC <= memory_to_writeBack_PC;
  writeBack_INSTRUCTION <= memory_to_writeBack_INSTRUCTION;
  process(when_DBusCachedPlugin_l307,switch_Fetcher_l362)
  begin
    decode_arbitration_haltItself <= pkg_toStdLogic(false);
    if when_DBusCachedPlugin_l307 = '1' then
      decode_arbitration_haltItself <= pkg_toStdLogic(true);
    end if;
    case switch_Fetcher_l362 is
      when "010" =>
        decode_arbitration_haltItself <= pkg_toStdLogic(true);
      when others =>
    end case;
  end process;

  process(when_HazardSimplePlugin_l113,CsrPlugin_pipelineLiberator_active,when_CsrPlugin_l1116)
  begin
    decode_arbitration_haltByOther <= pkg_toStdLogic(false);
    if when_HazardSimplePlugin_l113 = '1' then
      decode_arbitration_haltByOther <= pkg_toStdLogic(true);
    end if;
    if CsrPlugin_pipelineLiberator_active = '1' then
      decode_arbitration_haltByOther <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1116 = '1' then
      decode_arbitration_haltByOther <= pkg_toStdLogic(true);
    end if;
  end process;

  process(zz_when,decode_arbitration_isFlushed)
  begin
    decode_arbitration_removeIt <= pkg_toStdLogic(false);
    if zz_when = '1' then
      decode_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
    if decode_arbitration_isFlushed = '1' then
      decode_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
  end process;

  decode_arbitration_flushIt <= pkg_toStdLogic(false);
  process(zz_when)
  begin
    decode_arbitration_flushNext <= pkg_toStdLogic(false);
    if zz_when = '1' then
      decode_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DBusCachedPlugin_l347,when_CsrPlugin_l1180,execute_CsrPlugin_blockedBySideEffects)
  begin
    execute_arbitration_haltItself <= pkg_toStdLogic(false);
    if when_DBusCachedPlugin_l347 = '1' then
      execute_arbitration_haltItself <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1180 = '1' then
      if execute_CsrPlugin_blockedBySideEffects = '1' then
        execute_arbitration_haltItself <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  process(when_DBusCachedPlugin_l363,when_DebugPlugin_l295)
  begin
    execute_arbitration_haltByOther <= pkg_toStdLogic(false);
    if when_DBusCachedPlugin_l363 = '1' then
      execute_arbitration_haltByOther <= pkg_toStdLogic(true);
    end if;
    if when_DebugPlugin_l295 = '1' then
      execute_arbitration_haltByOther <= pkg_toStdLogic(true);
    end if;
  end process;

  process(execute_arbitration_isFlushed)
  begin
    execute_arbitration_removeIt <= pkg_toStdLogic(false);
    if execute_arbitration_isFlushed = '1' then
      execute_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DebugPlugin_l295,when_DebugPlugin_l298)
  begin
    execute_arbitration_flushIt <= pkg_toStdLogic(false);
    if when_DebugPlugin_l295 = '1' then
      if when_DebugPlugin_l298 = '1' then
        execute_arbitration_flushIt <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  process(when_DebugPlugin_l295,when_DebugPlugin_l298)
  begin
    execute_arbitration_flushNext <= pkg_toStdLogic(false);
    if when_DebugPlugin_l295 = '1' then
      if when_DebugPlugin_l298 = '1' then
        execute_arbitration_flushNext <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  process(when_MulDivIterativePlugin_l128,when_MulDivIterativePlugin_l129)
  begin
    memory_arbitration_haltItself <= pkg_toStdLogic(false);
    if when_MulDivIterativePlugin_l128 = '1' then
      if when_MulDivIterativePlugin_l129 = '1' then
        memory_arbitration_haltItself <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  memory_arbitration_haltByOther <= pkg_toStdLogic(false);
  process(BranchPlugin_branchExceptionPort_valid,memory_arbitration_isFlushed)
  begin
    memory_arbitration_removeIt <= pkg_toStdLogic(false);
    if BranchPlugin_branchExceptionPort_valid = '1' then
      memory_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
    if memory_arbitration_isFlushed = '1' then
      memory_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
  end process;

  memory_arbitration_flushIt <= pkg_toStdLogic(false);
  process(BranchPlugin_jumpInterface_valid,BranchPlugin_branchExceptionPort_valid)
  begin
    memory_arbitration_flushNext <= pkg_toStdLogic(false);
    if BranchPlugin_jumpInterface_valid = '1' then
      memory_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
    if BranchPlugin_branchExceptionPort_valid = '1' then
      memory_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DBusCachedPlugin_l462)
  begin
    writeBack_arbitration_haltItself <= pkg_toStdLogic(false);
    if when_DBusCachedPlugin_l462 = '1' then
      writeBack_arbitration_haltItself <= pkg_toStdLogic(true);
    end if;
  end process;

  writeBack_arbitration_haltByOther <= pkg_toStdLogic(false);
  process(DBusCachedPlugin_exceptionBus_valid,writeBack_arbitration_isFlushed)
  begin
    writeBack_arbitration_removeIt <= pkg_toStdLogic(false);
    if DBusCachedPlugin_exceptionBus_valid = '1' then
      writeBack_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
    if writeBack_arbitration_isFlushed = '1' then
      writeBack_arbitration_removeIt <= pkg_toStdLogic(true);
    end if;
  end process;

  process(DBusCachedPlugin_redoBranch_valid)
  begin
    writeBack_arbitration_flushIt <= pkg_toStdLogic(false);
    if DBusCachedPlugin_redoBranch_valid = '1' then
      writeBack_arbitration_flushIt <= pkg_toStdLogic(true);
    end if;
  end process;

  process(DBusCachedPlugin_redoBranch_valid,DBusCachedPlugin_exceptionBus_valid,when_CsrPlugin_l1019,when_CsrPlugin_l1064)
  begin
    writeBack_arbitration_flushNext <= pkg_toStdLogic(false);
    if DBusCachedPlugin_redoBranch_valid = '1' then
      writeBack_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
    if DBusCachedPlugin_exceptionBus_valid = '1' then
      writeBack_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1019 = '1' then
      writeBack_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1064 = '1' then
      writeBack_arbitration_flushNext <= pkg_toStdLogic(true);
    end if;
  end process;

  lastStageInstruction <= writeBack_INSTRUCTION;
  lastStagePc <= writeBack_PC;
  lastStageIsValid <= writeBack_arbitration_isValid;
  lastStageIsFiring <= writeBack_arbitration_isFiring;
  process(when_CsrPlugin_l922,when_CsrPlugin_l1019,when_CsrPlugin_l1064,when_DebugPlugin_l295,when_DebugPlugin_l298,DebugPlugin_haltIt,when_DebugPlugin_l311)
  begin
    IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(false);
    if when_CsrPlugin_l922 = '1' then
      IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1019 = '1' then
      IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1064 = '1' then
      IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(true);
    end if;
    if when_DebugPlugin_l295 = '1' then
      if when_DebugPlugin_l298 = '1' then
        IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(true);
      end if;
    end if;
    if DebugPlugin_haltIt = '1' then
      IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(true);
    end if;
    if when_DebugPlugin_l311 = '1' then
      IBusCachedPlugin_fetcherHalt <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_Fetcher_l240)
  begin
    IBusCachedPlugin_incomingInstruction <= pkg_toStdLogic(false);
    if when_Fetcher_l240 = '1' then
      IBusCachedPlugin_incomingInstruction <= pkg_toStdLogic(true);
    end if;
  end process;

  process(DebugPlugin_godmode)
  begin
    zz_when_DBusCachedPlugin_l390 <= pkg_toStdLogic(false);
    if DebugPlugin_godmode = '1' then
      zz_when_DBusCachedPlugin_l390 <= pkg_toStdLogic(true);
    end if;
  end process;

  CsrPlugin_csrMapping_allowCsrSignal <= pkg_toStdLogic(false);
  CsrPlugin_csrMapping_readDataSignal <= CsrPlugin_csrMapping_readDataInit;
  CsrPlugin_inWfi <= pkg_toStdLogic(false);
  process(DebugPlugin_haltIt)
  begin
    CsrPlugin_thirdPartyWake <= pkg_toStdLogic(false);
    if DebugPlugin_haltIt = '1' then
      CsrPlugin_thirdPartyWake <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_CsrPlugin_l1019,when_CsrPlugin_l1064)
  begin
    CsrPlugin_jumpInterface_valid <= pkg_toStdLogic(false);
    if when_CsrPlugin_l1019 = '1' then
      CsrPlugin_jumpInterface_valid <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1064 = '1' then
      CsrPlugin_jumpInterface_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_CsrPlugin_l1019,CsrPlugin_xtvec_base,when_CsrPlugin_l1064,switch_CsrPlugin_l1068,CsrPlugin_mepc)
  begin
    CsrPlugin_jumpInterface_payload <= pkg_unsigned("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
    if when_CsrPlugin_l1019 = '1' then
      CsrPlugin_jumpInterface_payload <= unsigned(pkg_cat(std_logic_vector(CsrPlugin_xtvec_base),std_logic_vector(pkg_unsigned("00"))));
    end if;
    if when_CsrPlugin_l1064 = '1' then
      case switch_CsrPlugin_l1068 is
        when "11" =>
          CsrPlugin_jumpInterface_payload <= CsrPlugin_mepc;
        when others =>
      end case;
    end if;
  end process;

  process(DebugPlugin_godmode)
  begin
    CsrPlugin_forceMachineWire <= pkg_toStdLogic(false);
    if DebugPlugin_godmode = '1' then
      CsrPlugin_forceMachineWire <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_DebugPlugin_l327)
  begin
    CsrPlugin_allowInterrupts <= pkg_toStdLogic(true);
    if when_DebugPlugin_l327 = '1' then
      CsrPlugin_allowInterrupts <= pkg_toStdLogic(false);
    end if;
  end process;

  process(DebugPlugin_godmode)
  begin
    CsrPlugin_allowException <= pkg_toStdLogic(true);
    if DebugPlugin_godmode = '1' then
      CsrPlugin_allowException <= pkg_toStdLogic(false);
    end if;
  end process;

  process(DebugPlugin_allowEBreak)
  begin
    CsrPlugin_allowEbreakException <= pkg_toStdLogic(true);
    if DebugPlugin_allowEBreak = '1' then
      CsrPlugin_allowEbreakException <= pkg_toStdLogic(false);
    end if;
  end process;

  IBusCachedPlugin_externalFlush <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_flushNext),pkg_cat(pkg_toStdLogicVector(memory_arbitration_flushNext),pkg_cat(pkg_toStdLogicVector(execute_arbitration_flushNext),pkg_toStdLogicVector(decode_arbitration_flushNext)))) /= pkg_stdLogicVector("0000"));
  IBusCachedPlugin_jump_pcLoad_valid <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(CsrPlugin_jumpInterface_valid),pkg_cat(pkg_toStdLogicVector(BranchPlugin_jumpInterface_valid),pkg_toStdLogicVector(DBusCachedPlugin_redoBranch_valid))) /= pkg_stdLogicVector("000"));
  zz_IBusCachedPlugin_jump_pcLoad_payload <= unsigned(pkg_cat(pkg_toStdLogicVector(BranchPlugin_jumpInterface_valid),pkg_cat(pkg_toStdLogicVector(CsrPlugin_jumpInterface_valid),pkg_toStdLogicVector(DBusCachedPlugin_redoBranch_valid))));
  zz_IBusCachedPlugin_jump_pcLoad_payload_1 <= std_logic_vector((zz_IBusCachedPlugin_jump_pcLoad_payload and pkg_not((zz_IBusCachedPlugin_jump_pcLoad_payload - pkg_unsigned("001")))));
  zz_IBusCachedPlugin_jump_pcLoad_payload_2 <= pkg_extract(zz_IBusCachedPlugin_jump_pcLoad_payload_1,1);
  zz_IBusCachedPlugin_jump_pcLoad_payload_3 <= pkg_extract(zz_IBusCachedPlugin_jump_pcLoad_payload_1,2);
  IBusCachedPlugin_jump_pcLoad_payload <= zz_IBusCachedPlugin_jump_pcLoad_payload_4;
  process(IBusCachedPlugin_fetchPc_predictionPcLoad_valid,IBusCachedPlugin_fetchPc_redo_valid,IBusCachedPlugin_jump_pcLoad_valid)
  begin
    IBusCachedPlugin_fetchPc_correction <= pkg_toStdLogic(false);
    if IBusCachedPlugin_fetchPc_predictionPcLoad_valid = '1' then
      IBusCachedPlugin_fetchPc_correction <= pkg_toStdLogic(true);
    end if;
    if IBusCachedPlugin_fetchPc_redo_valid = '1' then
      IBusCachedPlugin_fetchPc_correction <= pkg_toStdLogic(true);
    end if;
    if IBusCachedPlugin_jump_pcLoad_valid = '1' then
      IBusCachedPlugin_fetchPc_correction <= pkg_toStdLogic(true);
    end if;
  end process;

  IBusCachedPlugin_fetchPc_output_fire <= (IBusCachedPlugin_fetchPc_output_valid and IBusCachedPlugin_fetchPc_output_ready);
  IBusCachedPlugin_fetchPc_corrected <= (IBusCachedPlugin_fetchPc_correction or IBusCachedPlugin_fetchPc_correctionReg);
  IBusCachedPlugin_fetchPc_pcRegPropagate <= pkg_toStdLogic(false);
  when_Fetcher_l131 <= (IBusCachedPlugin_fetchPc_correction or IBusCachedPlugin_fetchPc_pcRegPropagate);
  IBusCachedPlugin_fetchPc_output_fire_1 <= (IBusCachedPlugin_fetchPc_output_valid and IBusCachedPlugin_fetchPc_output_ready);
  when_Fetcher_l131_1 <= ((not IBusCachedPlugin_fetchPc_output_valid) and IBusCachedPlugin_fetchPc_output_ready);
  process(IBusCachedPlugin_fetchPc_pcReg,IBusCachedPlugin_fetchPc_inc,IBusCachedPlugin_fetchPc_predictionPcLoad_valid,IBusCachedPlugin_fetchPc_predictionPcLoad_payload,IBusCachedPlugin_fetchPc_redo_valid,IBusCachedPlugin_fetchPc_redo_payload,IBusCachedPlugin_jump_pcLoad_valid,IBusCachedPlugin_jump_pcLoad_payload)
  begin
    IBusCachedPlugin_fetchPc_pc <= (IBusCachedPlugin_fetchPc_pcReg + pkg_resize(unsigned(pkg_cat(pkg_toStdLogicVector(IBusCachedPlugin_fetchPc_inc),pkg_stdLogicVector("00"))),32));
    if IBusCachedPlugin_fetchPc_predictionPcLoad_valid = '1' then
      IBusCachedPlugin_fetchPc_pc <= IBusCachedPlugin_fetchPc_predictionPcLoad_payload;
    end if;
    if IBusCachedPlugin_fetchPc_redo_valid = '1' then
      IBusCachedPlugin_fetchPc_pc <= IBusCachedPlugin_fetchPc_redo_payload;
    end if;
    if IBusCachedPlugin_jump_pcLoad_valid = '1' then
      IBusCachedPlugin_fetchPc_pc <= IBusCachedPlugin_jump_pcLoad_payload;
    end if;
    IBusCachedPlugin_fetchPc_pc(0) <= pkg_toStdLogic(false);
    IBusCachedPlugin_fetchPc_pc(1) <= pkg_toStdLogic(false);
  end process;

  process(IBusCachedPlugin_fetchPc_redo_valid,IBusCachedPlugin_jump_pcLoad_valid)
  begin
    IBusCachedPlugin_fetchPc_flushed <= pkg_toStdLogic(false);
    if IBusCachedPlugin_fetchPc_redo_valid = '1' then
      IBusCachedPlugin_fetchPc_flushed <= pkg_toStdLogic(true);
    end if;
    if IBusCachedPlugin_jump_pcLoad_valid = '1' then
      IBusCachedPlugin_fetchPc_flushed <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Fetcher_l158 <= (IBusCachedPlugin_fetchPc_booted and ((IBusCachedPlugin_fetchPc_output_ready or IBusCachedPlugin_fetchPc_correction) or IBusCachedPlugin_fetchPc_pcRegPropagate));
  IBusCachedPlugin_fetchPc_output_valid <= ((not IBusCachedPlugin_fetcherHalt) and IBusCachedPlugin_fetchPc_booted);
  IBusCachedPlugin_fetchPc_output_payload <= IBusCachedPlugin_fetchPc_pc;
  process(IBusCachedPlugin_rsp_redoFetch)
  begin
    IBusCachedPlugin_iBusRsp_redoFetch <= pkg_toStdLogic(false);
    if IBusCachedPlugin_rsp_redoFetch = '1' then
      IBusCachedPlugin_iBusRsp_redoFetch <= pkg_toStdLogic(true);
    end if;
  end process;

  IBusCachedPlugin_iBusRsp_stages_0_input_valid <= IBusCachedPlugin_fetchPc_output_valid;
  IBusCachedPlugin_fetchPc_output_ready <= IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  IBusCachedPlugin_iBusRsp_stages_0_input_payload <= IBusCachedPlugin_fetchPc_output_payload;
  process(IBusCachedPlugin_cache_io_cpu_prefetch_haltIt)
  begin
    IBusCachedPlugin_iBusRsp_stages_0_halt <= pkg_toStdLogic(false);
    if IBusCachedPlugin_cache_io_cpu_prefetch_haltIt = '1' then
      IBusCachedPlugin_iBusRsp_stages_0_halt <= pkg_toStdLogic(true);
    end if;
  end process;

  zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready <= (not IBusCachedPlugin_iBusRsp_stages_0_halt);
  IBusCachedPlugin_iBusRsp_stages_0_input_ready <= (IBusCachedPlugin_iBusRsp_stages_0_output_ready and zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  IBusCachedPlugin_iBusRsp_stages_0_output_valid <= (IBusCachedPlugin_iBusRsp_stages_0_input_valid and zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  IBusCachedPlugin_iBusRsp_stages_0_output_payload <= IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  process(IBusCachedPlugin_mmuBus_busy)
  begin
    IBusCachedPlugin_iBusRsp_stages_1_halt <= pkg_toStdLogic(false);
    if IBusCachedPlugin_mmuBus_busy = '1' then
      IBusCachedPlugin_iBusRsp_stages_1_halt <= pkg_toStdLogic(true);
    end if;
  end process;

  zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready <= (not IBusCachedPlugin_iBusRsp_stages_1_halt);
  IBusCachedPlugin_iBusRsp_stages_1_input_ready <= (IBusCachedPlugin_iBusRsp_stages_1_output_ready and zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  IBusCachedPlugin_iBusRsp_stages_1_output_valid <= (IBusCachedPlugin_iBusRsp_stages_1_input_valid and zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  IBusCachedPlugin_iBusRsp_stages_1_output_payload <= IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  process(when_IBusCachedPlugin_l267)
  begin
    IBusCachedPlugin_iBusRsp_stages_2_halt <= pkg_toStdLogic(false);
    if when_IBusCachedPlugin_l267 = '1' then
      IBusCachedPlugin_iBusRsp_stages_2_halt <= pkg_toStdLogic(true);
    end if;
  end process;

  zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready <= (not IBusCachedPlugin_iBusRsp_stages_2_halt);
  IBusCachedPlugin_iBusRsp_stages_2_input_ready <= (IBusCachedPlugin_iBusRsp_stages_2_output_ready and zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  IBusCachedPlugin_iBusRsp_stages_2_output_valid <= (IBusCachedPlugin_iBusRsp_stages_2_input_valid and zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  IBusCachedPlugin_iBusRsp_stages_2_output_payload <= IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  IBusCachedPlugin_fetchPc_redo_valid <= IBusCachedPlugin_iBusRsp_redoFetch;
  IBusCachedPlugin_fetchPc_redo_payload <= IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  IBusCachedPlugin_iBusRsp_flush <= ((decode_arbitration_removeIt or (decode_arbitration_flushNext and (not decode_arbitration_isStuck))) or IBusCachedPlugin_iBusRsp_redoFetch);
  IBusCachedPlugin_iBusRsp_stages_0_output_ready <= ((pkg_toStdLogic(false) and (not IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid)) or IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_ready);
  IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid <= zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid;
  IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_payload <= zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_payload;
  IBusCachedPlugin_iBusRsp_stages_1_input_valid <= IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid;
  IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_ready <= IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  IBusCachedPlugin_iBusRsp_stages_1_input_payload <= IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_payload;
  IBusCachedPlugin_iBusRsp_stages_1_output_ready <= ((pkg_toStdLogic(false) and (not IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid)) or IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready);
  IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  IBusCachedPlugin_iBusRsp_stages_2_input_valid <= IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready <= IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  IBusCachedPlugin_iBusRsp_stages_2_input_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  process(when_Fetcher_l320)
  begin
    IBusCachedPlugin_iBusRsp_readyForError <= pkg_toStdLogic(true);
    if when_Fetcher_l320 = '1' then
      IBusCachedPlugin_iBusRsp_readyForError <= pkg_toStdLogic(false);
    end if;
  end process;

  when_Fetcher_l240 <= (IBusCachedPlugin_iBusRsp_stages_1_input_valid or IBusCachedPlugin_iBusRsp_stages_2_input_valid);
  when_Fetcher_l320 <= (not IBusCachedPlugin_pcValids_0);
  when_Fetcher_l329 <= (not (not IBusCachedPlugin_iBusRsp_stages_1_input_ready));
  when_Fetcher_l329_1 <= (not (not IBusCachedPlugin_iBusRsp_stages_2_input_ready));
  when_Fetcher_l329_2 <= (not execute_arbitration_isStuck);
  when_Fetcher_l329_3 <= (not memory_arbitration_isStuck);
  when_Fetcher_l329_4 <= (not writeBack_arbitration_isStuck);
  IBusCachedPlugin_pcValids_0 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
  IBusCachedPlugin_pcValids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
  IBusCachedPlugin_pcValids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_3;
  IBusCachedPlugin_pcValids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_4;
  IBusCachedPlugin_iBusRsp_output_ready <= (not decode_arbitration_isStuck);
  process(IBusCachedPlugin_iBusRsp_output_valid,switch_Fetcher_l362)
  begin
    decode_arbitration_isValid <= IBusCachedPlugin_iBusRsp_output_valid;
    case switch_Fetcher_l362 is
      when "010" =>
        decode_arbitration_isValid <= pkg_toStdLogic(true);
      when "011" =>
        decode_arbitration_isValid <= pkg_toStdLogic(true);
      when others =>
    end case;
  end process;

  IBusCachedPlugin_predictor_historyWriteDelayPatched_valid <= IBusCachedPlugin_predictor_historyWrite_valid;
  IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_address <= (IBusCachedPlugin_predictor_historyWrite_payload_address - pkg_unsigned("00000001"));
  IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_source <= IBusCachedPlugin_predictor_historyWrite_payload_data_source;
  IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_branchWish <= IBusCachedPlugin_predictor_historyWrite_payload_data_branchWish;
  IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_target <= IBusCachedPlugin_predictor_historyWrite_payload_data_target;
  zz_IBusCachedPlugin_predictor_buffer_line_source <= pkg_shiftRight(IBusCachedPlugin_iBusRsp_stages_0_input_payload,2);
  zz_IBusCachedPlugin_predictor_buffer_line_source_1 <= zz_IBusCachedPlugin_predictor_history_port0;
  IBusCachedPlugin_predictor_buffer_line_source <= pkg_extract(zz_IBusCachedPlugin_predictor_buffer_line_source_1,21,0);
  IBusCachedPlugin_predictor_buffer_line_branchWish <= unsigned(pkg_extract(zz_IBusCachedPlugin_predictor_buffer_line_source_1,23,22));
  IBusCachedPlugin_predictor_buffer_line_target <= unsigned(pkg_extract(zz_IBusCachedPlugin_predictor_buffer_line_source_1,55,24));
  IBusCachedPlugin_predictor_buffer_hazard <= (IBusCachedPlugin_predictor_writeLast_valid and pkg_toStdLogic(IBusCachedPlugin_predictor_writeLast_payload_address = pkg_resize(pkg_shiftRight(IBusCachedPlugin_iBusRsp_stages_1_input_payload,2),8)));
  IBusCachedPlugin_predictor_hazard <= (IBusCachedPlugin_predictor_buffer_hazard_regNextWhen or IBusCachedPlugin_predictor_buffer_pcCorrected);
  IBusCachedPlugin_predictor_hit <= pkg_toStdLogic(IBusCachedPlugin_predictor_line_source = pkg_shiftRight(std_logic_vector(IBusCachedPlugin_iBusRsp_stages_1_input_payload),10));
  IBusCachedPlugin_fetchPc_predictionPcLoad_valid <= (((pkg_extract(IBusCachedPlugin_predictor_line_branchWish,1) and IBusCachedPlugin_predictor_hit) and (not IBusCachedPlugin_predictor_hazard)) and IBusCachedPlugin_iBusRsp_stages_1_input_valid);
  IBusCachedPlugin_fetchPc_predictionPcLoad_payload <= IBusCachedPlugin_predictor_line_target;
  IBusCachedPlugin_predictor_fetchContext_hazard <= IBusCachedPlugin_predictor_hazard;
  IBusCachedPlugin_predictor_fetchContext_hit <= IBusCachedPlugin_predictor_hit;
  IBusCachedPlugin_predictor_fetchContext_line_source <= IBusCachedPlugin_predictor_line_source;
  IBusCachedPlugin_predictor_fetchContext_line_branchWish <= IBusCachedPlugin_predictor_line_branchWish;
  IBusCachedPlugin_predictor_fetchContext_line_target <= IBusCachedPlugin_predictor_line_target;
  IBusCachedPlugin_predictor_iBusRspContextOutput_hazard <= IBusCachedPlugin_predictor_iBusRspContext_hazard;
  IBusCachedPlugin_predictor_iBusRspContextOutput_hit <= IBusCachedPlugin_predictor_iBusRspContext_hit;
  IBusCachedPlugin_predictor_iBusRspContextOutput_line_source <= IBusCachedPlugin_predictor_iBusRspContext_line_source;
  IBusCachedPlugin_predictor_iBusRspContextOutput_line_branchWish <= IBusCachedPlugin_predictor_iBusRspContext_line_branchWish;
  IBusCachedPlugin_predictor_iBusRspContextOutput_line_target <= IBusCachedPlugin_predictor_iBusRspContext_line_target;
  IBusCachedPlugin_predictor_injectorContext_hazard <= IBusCachedPlugin_predictor_iBusRspContextOutput_hazard;
  IBusCachedPlugin_predictor_injectorContext_hit <= IBusCachedPlugin_predictor_iBusRspContextOutput_hit;
  IBusCachedPlugin_predictor_injectorContext_line_source <= IBusCachedPlugin_predictor_iBusRspContextOutput_line_source;
  IBusCachedPlugin_predictor_injectorContext_line_branchWish <= IBusCachedPlugin_predictor_iBusRspContextOutput_line_branchWish;
  IBusCachedPlugin_predictor_injectorContext_line_target <= IBusCachedPlugin_predictor_iBusRspContextOutput_line_target;
  IBusCachedPlugin_fetchPrediction_cmd_hadBranch <= ((memory_PREDICTION_CONTEXT_hit and (not memory_PREDICTION_CONTEXT_hazard)) and pkg_extract(memory_PREDICTION_CONTEXT_line_branchWish,1));
  IBusCachedPlugin_fetchPrediction_cmd_targetPc <= memory_PREDICTION_CONTEXT_line_target;
  process(IBusCachedPlugin_fetchPrediction_rsp_wasRight,memory_PREDICTION_CONTEXT_hit,when_Fetcher_l596)
  begin
    IBusCachedPlugin_predictor_historyWrite_valid <= pkg_toStdLogic(false);
    if IBusCachedPlugin_fetchPrediction_rsp_wasRight = '1' then
      IBusCachedPlugin_predictor_historyWrite_valid <= memory_PREDICTION_CONTEXT_hit;
    else
      if memory_PREDICTION_CONTEXT_hit = '1' then
        IBusCachedPlugin_predictor_historyWrite_valid <= pkg_toStdLogic(true);
      else
        IBusCachedPlugin_predictor_historyWrite_valid <= pkg_toStdLogic(true);
      end if;
    end if;
    if when_Fetcher_l596 = '1' then
      IBusCachedPlugin_predictor_historyWrite_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  IBusCachedPlugin_predictor_historyWrite_payload_address <= pkg_extract(IBusCachedPlugin_fetchPrediction_rsp_sourceLastWord,9,2);
  IBusCachedPlugin_predictor_historyWrite_payload_data_source <= pkg_shiftRight(std_logic_vector(IBusCachedPlugin_fetchPrediction_rsp_sourceLastWord),10);
  IBusCachedPlugin_predictor_historyWrite_payload_data_target <= IBusCachedPlugin_fetchPrediction_rsp_finalPc;
  process(IBusCachedPlugin_fetchPrediction_rsp_wasRight,memory_PREDICTION_CONTEXT_line_branchWish,memory_PREDICTION_CONTEXT_hit)
  begin
    if IBusCachedPlugin_fetchPrediction_rsp_wasRight = '1' then
      IBusCachedPlugin_predictor_historyWrite_payload_data_branchWish <= ((memory_PREDICTION_CONTEXT_line_branchWish + pkg_resize(unsigned(pkg_toStdLogicVector(pkg_toStdLogic(memory_PREDICTION_CONTEXT_line_branchWish = pkg_unsigned("10")))),2)) - pkg_resize(unsigned(pkg_toStdLogicVector(pkg_toStdLogic(memory_PREDICTION_CONTEXT_line_branchWish = pkg_unsigned("01")))),2));
    else
      if memory_PREDICTION_CONTEXT_hit = '1' then
        IBusCachedPlugin_predictor_historyWrite_payload_data_branchWish <= ((memory_PREDICTION_CONTEXT_line_branchWish - pkg_resize(unsigned(pkg_toStdLogicVector(pkg_extract(memory_PREDICTION_CONTEXT_line_branchWish,1))),2)) + pkg_resize(unsigned(pkg_toStdLogicVector((not pkg_extract(memory_PREDICTION_CONTEXT_line_branchWish,1)))),2));
      else
        IBusCachedPlugin_predictor_historyWrite_payload_data_branchWish <= pkg_unsigned("10");
      end if;
    end if;
  end process;

  when_Fetcher_l596 <= (memory_PREDICTION_CONTEXT_hazard or (not memory_arbitration_isFiring));
  iBus_cmd_valid <= IBusCachedPlugin_cache_io_mem_cmd_valid;
  process(IBusCachedPlugin_cache_io_mem_cmd_payload_address)
  begin
    iBus_cmd_payload_address <= IBusCachedPlugin_cache_io_mem_cmd_payload_address;
    iBus_cmd_payload_address <= IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  end process;

  iBus_cmd_payload_size <= IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  IBusCachedPlugin_s0_tightlyCoupledHit <= pkg_toStdLogic(false);
  IBusCachedPlugin_cache_io_cpu_prefetch_isValid <= (IBusCachedPlugin_iBusRsp_stages_0_input_valid and (not IBusCachedPlugin_s0_tightlyCoupledHit));
  IBusCachedPlugin_cache_io_cpu_fetch_isValid <= (IBusCachedPlugin_iBusRsp_stages_1_input_valid and (not IBusCachedPlugin_s1_tightlyCoupledHit));
  IBusCachedPlugin_cache_io_cpu_fetch_isStuck <= (not IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  IBusCachedPlugin_mmuBus_cmd_0_isValid <= IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  IBusCachedPlugin_mmuBus_cmd_0_isStuck <= (not IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  IBusCachedPlugin_mmuBus_cmd_0_virtualAddress <= IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation <= pkg_toStdLogic(false);
  IBusCachedPlugin_mmuBus_end <= (IBusCachedPlugin_iBusRsp_stages_1_input_ready or IBusCachedPlugin_externalFlush);
  IBusCachedPlugin_cache_io_cpu_decode_isValid <= (IBusCachedPlugin_iBusRsp_stages_2_input_valid and (not IBusCachedPlugin_s2_tightlyCoupledHit));
  IBusCachedPlugin_cache_io_cpu_decode_isStuck <= (not IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  IBusCachedPlugin_cache_io_cpu_decode_isUser <= pkg_toStdLogic(CsrPlugin_privilege = pkg_unsigned("00"));
  IBusCachedPlugin_rsp_iBusRspOutputHalt <= pkg_toStdLogic(false);
  IBusCachedPlugin_rsp_issueDetected <= pkg_toStdLogic(false);
  process(when_IBusCachedPlugin_l239,when_IBusCachedPlugin_l250)
  begin
    IBusCachedPlugin_rsp_redoFetch <= pkg_toStdLogic(false);
    if when_IBusCachedPlugin_l239 = '1' then
      IBusCachedPlugin_rsp_redoFetch <= pkg_toStdLogic(true);
    end if;
    if when_IBusCachedPlugin_l250 = '1' then
      IBusCachedPlugin_rsp_redoFetch <= pkg_toStdLogic(true);
    end if;
  end process;

  process(IBusCachedPlugin_rsp_redoFetch,IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling,when_IBusCachedPlugin_l250)
  begin
    IBusCachedPlugin_cache_io_cpu_fill_valid <= (IBusCachedPlugin_rsp_redoFetch and (not IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling));
    if when_IBusCachedPlugin_l250 = '1' then
      IBusCachedPlugin_cache_io_cpu_fill_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_IBusCachedPlugin_l244,IBusCachedPlugin_iBusRsp_readyForError,when_IBusCachedPlugin_l256)
  begin
    IBusCachedPlugin_decodeExceptionPort_valid <= pkg_toStdLogic(false);
    if when_IBusCachedPlugin_l244 = '1' then
      IBusCachedPlugin_decodeExceptionPort_valid <= IBusCachedPlugin_iBusRsp_readyForError;
    end if;
    if when_IBusCachedPlugin_l256 = '1' then
      IBusCachedPlugin_decodeExceptionPort_valid <= IBusCachedPlugin_iBusRsp_readyForError;
    end if;
  end process;

  process(when_IBusCachedPlugin_l244,when_IBusCachedPlugin_l256)
  begin
    IBusCachedPlugin_decodeExceptionPort_payload_code <= pkg_unsigned("XXXX");
    if when_IBusCachedPlugin_l244 = '1' then
      IBusCachedPlugin_decodeExceptionPort_payload_code <= pkg_unsigned("1100");
    end if;
    if when_IBusCachedPlugin_l256 = '1' then
      IBusCachedPlugin_decodeExceptionPort_payload_code <= pkg_unsigned("0001");
    end if;
  end process;

  IBusCachedPlugin_decodeExceptionPort_payload_badAddr <= unsigned(pkg_cat(std_logic_vector(pkg_extract(IBusCachedPlugin_iBusRsp_stages_2_input_payload,31,2)),std_logic_vector(pkg_unsigned("00"))));
  when_IBusCachedPlugin_l239 <= ((IBusCachedPlugin_cache_io_cpu_decode_isValid and IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling) and (not IBusCachedPlugin_rsp_issueDetected));
  when_IBusCachedPlugin_l244 <= ((IBusCachedPlugin_cache_io_cpu_decode_isValid and IBusCachedPlugin_cache_io_cpu_decode_mmuException) and (not IBusCachedPlugin_rsp_issueDetected_1));
  when_IBusCachedPlugin_l250 <= ((IBusCachedPlugin_cache_io_cpu_decode_isValid and IBusCachedPlugin_cache_io_cpu_decode_cacheMiss) and (not IBusCachedPlugin_rsp_issueDetected_2));
  when_IBusCachedPlugin_l256 <= ((IBusCachedPlugin_cache_io_cpu_decode_isValid and IBusCachedPlugin_cache_io_cpu_decode_error) and (not IBusCachedPlugin_rsp_issueDetected_3));
  when_IBusCachedPlugin_l267 <= (IBusCachedPlugin_rsp_issueDetected_4 or IBusCachedPlugin_rsp_iBusRspOutputHalt);
  IBusCachedPlugin_iBusRsp_output_valid <= IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  IBusCachedPlugin_iBusRsp_stages_2_output_ready <= IBusCachedPlugin_iBusRsp_output_ready;
  IBusCachedPlugin_iBusRsp_output_payload_rsp_inst <= IBusCachedPlugin_cache_io_cpu_decode_data;
  IBusCachedPlugin_iBusRsp_output_payload_pc <= IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  IBusCachedPlugin_cache_io_flush <= (decode_arbitration_isValid and decode_FLUSH_ALL);
  dBus_cmd_valid <= dataCache_1_io_mem_cmd_valid;
  dBus_cmd_payload_wr <= dataCache_1_io_mem_cmd_payload_wr;
  dBus_cmd_payload_uncached <= dataCache_1_io_mem_cmd_payload_uncached;
  dBus_cmd_payload_address <= dataCache_1_io_mem_cmd_payload_address;
  dBus_cmd_payload_data <= dataCache_1_io_mem_cmd_payload_data;
  dBus_cmd_payload_mask <= dataCache_1_io_mem_cmd_payload_mask;
  dBus_cmd_payload_size <= dataCache_1_io_mem_cmd_payload_size;
  dBus_cmd_payload_last <= dataCache_1_io_mem_cmd_payload_last;
  when_DBusCachedPlugin_l307 <= ((DBusCachedPlugin_mmuBus_busy and decode_arbitration_isValid) and decode_MEMORY_ENABLE);
  execute_DBusCachedPlugin_size <= unsigned(pkg_extract(execute_INSTRUCTION,13,12));
  dataCache_1_io_cpu_execute_isValid <= (execute_arbitration_isValid and execute_MEMORY_ENABLE);
  dataCache_1_io_cpu_execute_address <= unsigned(execute_SRC_ADD);
  process(execute_DBusCachedPlugin_size,execute_RS2)
  begin
    case execute_DBusCachedPlugin_size is
      when "00" =>
        zz_execute_MEMORY_STORE_DATA_RF <= pkg_cat(pkg_cat(pkg_cat(pkg_extract(execute_RS2,7,0),pkg_extract(execute_RS2,7,0)),pkg_extract(execute_RS2,7,0)),pkg_extract(execute_RS2,7,0));
      when "01" =>
        zz_execute_MEMORY_STORE_DATA_RF <= pkg_cat(pkg_extract(execute_RS2,15,0),pkg_extract(execute_RS2,15,0));
      when others =>
        zz_execute_MEMORY_STORE_DATA_RF <= pkg_extract(execute_RS2,31,0);
    end case;
  end process;

  dataCache_1_io_cpu_flush_valid <= (execute_arbitration_isValid and execute_MEMORY_MANAGMENT);
  dataCache_1_io_cpu_flush_isStall <= (dataCache_1_io_cpu_flush_valid and (not dataCache_1_io_cpu_flush_ready));
  when_DBusCachedPlugin_l347 <= (dataCache_1_io_cpu_flush_isStall or dataCache_1_io_cpu_execute_haltIt);
  when_DBusCachedPlugin_l363 <= (dataCache_1_io_cpu_execute_refilling and execute_arbitration_isValid);
  dataCache_1_io_cpu_memory_isValid <= (memory_arbitration_isValid and memory_MEMORY_ENABLE);
  dataCache_1_io_cpu_memory_address <= unsigned(memory_REGFILE_WRITE_DATA);
  DBusCachedPlugin_mmuBus_cmd_0_isValid <= dataCache_1_io_cpu_memory_isValid;
  DBusCachedPlugin_mmuBus_cmd_0_isStuck <= memory_arbitration_isStuck;
  DBusCachedPlugin_mmuBus_cmd_0_virtualAddress <= dataCache_1_io_cpu_memory_address;
  DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation <= pkg_toStdLogic(false);
  DBusCachedPlugin_mmuBus_end <= ((not memory_arbitration_isStuck) or memory_arbitration_removeIt);
  process(DBusCachedPlugin_mmuBus_rsp_isIoAccess,when_DBusCachedPlugin_l390)
  begin
    dataCache_1_io_cpu_memory_mmuRsp_isIoAccess <= DBusCachedPlugin_mmuBus_rsp_isIoAccess;
    if when_DBusCachedPlugin_l390 = '1' then
      dataCache_1_io_cpu_memory_mmuRsp_isIoAccess <= pkg_toStdLogic(true);
    end if;
  end process;

  when_DBusCachedPlugin_l390 <= (zz_when_DBusCachedPlugin_l390 and (not dataCache_1_io_cpu_memory_isWrite));
  process(writeBack_arbitration_isValid,writeBack_MEMORY_ENABLE,writeBack_arbitration_haltByOther)
  begin
    dataCache_1_io_cpu_writeBack_isValid <= (writeBack_arbitration_isValid and writeBack_MEMORY_ENABLE);
    if writeBack_arbitration_haltByOther = '1' then
      dataCache_1_io_cpu_writeBack_isValid <= pkg_toStdLogic(false);
    end if;
  end process;

  dataCache_1_io_cpu_writeBack_isUser <= pkg_toStdLogic(CsrPlugin_privilege = pkg_unsigned("00"));
  dataCache_1_io_cpu_writeBack_address <= unsigned(writeBack_REGFILE_WRITE_DATA);
  dataCache_1_io_cpu_writeBack_storeData(31 downto 0) <= writeBack_MEMORY_STORE_DATA_RF;
  process(when_DBusCachedPlugin_l442,dataCache_1_io_cpu_redo)
  begin
    DBusCachedPlugin_redoBranch_valid <= pkg_toStdLogic(false);
    if when_DBusCachedPlugin_l442 = '1' then
      if dataCache_1_io_cpu_redo = '1' then
        DBusCachedPlugin_redoBranch_valid <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  DBusCachedPlugin_redoBranch_payload <= writeBack_PC;
  process(when_DBusCachedPlugin_l442,dataCache_1_io_cpu_writeBack_accessError,dataCache_1_io_cpu_writeBack_mmuException,dataCache_1_io_cpu_writeBack_unalignedAccess,dataCache_1_io_cpu_redo)
  begin
    DBusCachedPlugin_exceptionBus_valid <= pkg_toStdLogic(false);
    if when_DBusCachedPlugin_l442 = '1' then
      if dataCache_1_io_cpu_writeBack_accessError = '1' then
        DBusCachedPlugin_exceptionBus_valid <= pkg_toStdLogic(true);
      end if;
      if dataCache_1_io_cpu_writeBack_mmuException = '1' then
        DBusCachedPlugin_exceptionBus_valid <= pkg_toStdLogic(true);
      end if;
      if dataCache_1_io_cpu_writeBack_unalignedAccess = '1' then
        DBusCachedPlugin_exceptionBus_valid <= pkg_toStdLogic(true);
      end if;
      if dataCache_1_io_cpu_redo = '1' then
        DBusCachedPlugin_exceptionBus_valid <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

  DBusCachedPlugin_exceptionBus_payload_badAddr <= unsigned(writeBack_REGFILE_WRITE_DATA);
  process(when_DBusCachedPlugin_l442,dataCache_1_io_cpu_writeBack_accessError,writeBack_MEMORY_WR,dataCache_1_io_cpu_writeBack_mmuException,dataCache_1_io_cpu_writeBack_unalignedAccess)
  begin
    DBusCachedPlugin_exceptionBus_payload_code <= pkg_unsigned("XXXX");
    if when_DBusCachedPlugin_l442 = '1' then
      if dataCache_1_io_cpu_writeBack_accessError = '1' then
        DBusCachedPlugin_exceptionBus_payload_code <= pkg_resize(pkg_mux(writeBack_MEMORY_WR,pkg_unsigned("111"),pkg_unsigned("101")),4);
      end if;
      if dataCache_1_io_cpu_writeBack_mmuException = '1' then
        DBusCachedPlugin_exceptionBus_payload_code <= pkg_mux(writeBack_MEMORY_WR,pkg_unsigned("1111"),pkg_unsigned("1101"));
      end if;
      if dataCache_1_io_cpu_writeBack_unalignedAccess = '1' then
        DBusCachedPlugin_exceptionBus_payload_code <= pkg_resize(pkg_mux(writeBack_MEMORY_WR,pkg_unsigned("110"),pkg_unsigned("100")),4);
      end if;
    end if;
  end process;

  when_DBusCachedPlugin_l442 <= (writeBack_arbitration_isValid and writeBack_MEMORY_ENABLE);
  when_DBusCachedPlugin_l462 <= (dataCache_1_io_cpu_writeBack_isValid and dataCache_1_io_cpu_writeBack_haltIt);
  writeBack_DBusCachedPlugin_rspSplits_0 <= pkg_extract(dataCache_1_io_cpu_writeBack_data,7,0);
  writeBack_DBusCachedPlugin_rspSplits_1 <= pkg_extract(dataCache_1_io_cpu_writeBack_data,15,8);
  writeBack_DBusCachedPlugin_rspSplits_2 <= pkg_extract(dataCache_1_io_cpu_writeBack_data,23,16);
  writeBack_DBusCachedPlugin_rspSplits_3 <= pkg_extract(dataCache_1_io_cpu_writeBack_data,31,24);
  process(zz_writeBack_DBusCachedPlugin_rspShifted,zz_writeBack_DBusCachedPlugin_rspShifted_2,writeBack_DBusCachedPlugin_rspSplits_2,writeBack_DBusCachedPlugin_rspSplits_3)
  begin
    writeBack_DBusCachedPlugin_rspShifted(7 downto 0) <= zz_writeBack_DBusCachedPlugin_rspShifted;
    writeBack_DBusCachedPlugin_rspShifted(15 downto 8) <= zz_writeBack_DBusCachedPlugin_rspShifted_2;
    writeBack_DBusCachedPlugin_rspShifted(23 downto 16) <= writeBack_DBusCachedPlugin_rspSplits_2;
    writeBack_DBusCachedPlugin_rspShifted(31 downto 24) <= writeBack_DBusCachedPlugin_rspSplits_3;
  end process;

  writeBack_DBusCachedPlugin_rspRf <= pkg_extract(writeBack_DBusCachedPlugin_rspShifted,31,0);
  switch_Misc_l204 <= pkg_extract(writeBack_INSTRUCTION,13,12);
  zz_writeBack_DBusCachedPlugin_rspFormated <= (pkg_extract(writeBack_DBusCachedPlugin_rspRf,7) and (not pkg_extract(writeBack_INSTRUCTION,14)));
  process(zz_writeBack_DBusCachedPlugin_rspFormated,writeBack_DBusCachedPlugin_rspRf)
  begin
    zz_writeBack_DBusCachedPlugin_rspFormated_1(31) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(30) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(29) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(28) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(27) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(26) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(25) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(24) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(23) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(22) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(21) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(20) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(19) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(18) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(17) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(16) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(15) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(14) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(13) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(12) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(11) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(10) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(9) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(8) <= zz_writeBack_DBusCachedPlugin_rspFormated;
    zz_writeBack_DBusCachedPlugin_rspFormated_1(7 downto 0) <= pkg_extract(writeBack_DBusCachedPlugin_rspRf,7,0);
  end process;

  zz_writeBack_DBusCachedPlugin_rspFormated_2 <= (pkg_extract(writeBack_DBusCachedPlugin_rspRf,15) and (not pkg_extract(writeBack_INSTRUCTION,14)));
  process(zz_writeBack_DBusCachedPlugin_rspFormated_2,writeBack_DBusCachedPlugin_rspRf)
  begin
    zz_writeBack_DBusCachedPlugin_rspFormated_3(31) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(30) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(29) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(28) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(27) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(26) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(25) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(24) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(23) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(22) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(21) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(20) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(19) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(18) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(17) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(16) <= zz_writeBack_DBusCachedPlugin_rspFormated_2;
    zz_writeBack_DBusCachedPlugin_rspFormated_3(15 downto 0) <= pkg_extract(writeBack_DBusCachedPlugin_rspRf,15,0);
  end process;

  process(switch_Misc_l204,zz_writeBack_DBusCachedPlugin_rspFormated_1,zz_writeBack_DBusCachedPlugin_rspFormated_3,writeBack_DBusCachedPlugin_rspRf)
  begin
    case switch_Misc_l204 is
      when "00" =>
        writeBack_DBusCachedPlugin_rspFormated <= zz_writeBack_DBusCachedPlugin_rspFormated_1;
      when "01" =>
        writeBack_DBusCachedPlugin_rspFormated <= zz_writeBack_DBusCachedPlugin_rspFormated_3;
      when others =>
        writeBack_DBusCachedPlugin_rspFormated <= writeBack_DBusCachedPlugin_rspRf;
    end case;
  end process;

  when_DBusCachedPlugin_l488 <= (writeBack_arbitration_isValid and writeBack_MEMORY_ENABLE);
  IBusCachedPlugin_mmuBus_rsp_physicalAddress <= IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  IBusCachedPlugin_mmuBus_rsp_allowRead <= pkg_toStdLogic(true);
  IBusCachedPlugin_mmuBus_rsp_allowWrite <= pkg_toStdLogic(true);
  IBusCachedPlugin_mmuBus_rsp_allowExecute <= pkg_toStdLogic(true);
  IBusCachedPlugin_mmuBus_rsp_isIoAccess <= pkg_toStdLogic(pkg_extract(IBusCachedPlugin_mmuBus_rsp_physicalAddress,31,28) = pkg_unsigned("1111"));
  IBusCachedPlugin_mmuBus_rsp_isPaging <= pkg_toStdLogic(false);
  IBusCachedPlugin_mmuBus_rsp_exception <= pkg_toStdLogic(false);
  IBusCachedPlugin_mmuBus_rsp_refilling <= pkg_toStdLogic(false);
  IBusCachedPlugin_mmuBus_busy <= pkg_toStdLogic(false);
  DBusCachedPlugin_mmuBus_rsp_physicalAddress <= DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  DBusCachedPlugin_mmuBus_rsp_allowRead <= pkg_toStdLogic(true);
  DBusCachedPlugin_mmuBus_rsp_allowWrite <= pkg_toStdLogic(true);
  DBusCachedPlugin_mmuBus_rsp_allowExecute <= pkg_toStdLogic(true);
  DBusCachedPlugin_mmuBus_rsp_isIoAccess <= pkg_toStdLogic(pkg_extract(DBusCachedPlugin_mmuBus_rsp_physicalAddress,31,28) = pkg_unsigned("1111"));
  DBusCachedPlugin_mmuBus_rsp_isPaging <= pkg_toStdLogic(false);
  DBusCachedPlugin_mmuBus_rsp_exception <= pkg_toStdLogic(false);
  DBusCachedPlugin_mmuBus_rsp_refilling <= pkg_toStdLogic(false);
  DBusCachedPlugin_mmuBus_busy <= pkg_toStdLogic(false);
  zz_decode_ENV_CTRL_3 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000100000001010000")) = pkg_stdLogicVector("00000000000000000100000001010000"));
  zz_decode_ENV_CTRL_4 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000011000")) = pkg_stdLogicVector("00000000000000000000000000000000"));
  zz_decode_ENV_CTRL_5 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000000100")) = pkg_stdLogicVector("00000000000000000000000000000100"));
  zz_decode_ENV_CTRL_6 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000001001000")) = pkg_stdLogicVector("00000000000000000000000001001000"));
  zz_decode_ENV_CTRL_7 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000000000000110000")) = pkg_stdLogicVector("00000000000000000000000000010000"));
  zz_decode_ENV_CTRL_8 <= pkg_toStdLogic((decode_INSTRUCTION and pkg_stdLogicVector("00000000000000000001000000000000")) = pkg_stdLogicVector("00000000000000000000000000000000"));
  zz_decode_ENV_CTRL_2 <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic((decode_INSTRUCTION and zz_zz_decode_ENV_CTRL_2) = pkg_stdLogicVector("00000000000000000000000001010000"))) /= pkg_stdLogicVector("0"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_1 = zz_zz_decode_ENV_CTRL_2_2)) /= pkg_stdLogicVector("0"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(pkg_cat(zz_zz_decode_ENV_CTRL_2_3,zz_zz_decode_ENV_CTRL_2_5) /= pkg_stdLogicVector("00"))),pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(zz_zz_decode_ENV_CTRL_2_7 /= zz_zz_decode_ENV_CTRL_2_10)),pkg_cat(pkg_toStdLogicVector(zz_zz_decode_ENV_CTRL_2_11),pkg_cat(zz_zz_decode_ENV_CTRL_2_14,zz_zz_decode_ENV_CTRL_2_15))))));
  zz_decode_SRC1_CTRL_2 <= pkg_extract(zz_decode_ENV_CTRL_2,2,1);
  zz_decode_SRC1_CTRL_1 <= zz_decode_SRC1_CTRL_2;
  zz_decode_ALU_CTRL_2 <= pkg_extract(zz_decode_ENV_CTRL_2,7,6);
  zz_decode_ALU_CTRL_1 <= zz_decode_ALU_CTRL_2;
  zz_decode_SRC2_CTRL_2 <= pkg_extract(zz_decode_ENV_CTRL_2,9,8);
  zz_decode_SRC2_CTRL_1 <= zz_decode_SRC2_CTRL_2;
  zz_decode_ALU_BITWISE_CTRL_2 <= pkg_extract(zz_decode_ENV_CTRL_2,19,18);
  zz_decode_ALU_BITWISE_CTRL_1 <= zz_decode_ALU_BITWISE_CTRL_2;
  zz_decode_SHIFT_CTRL_2 <= pkg_extract(zz_decode_ENV_CTRL_2,22,21);
  zz_decode_SHIFT_CTRL_1 <= zz_decode_SHIFT_CTRL_2;
  zz_decode_BRANCH_CTRL_2 <= pkg_extract(zz_decode_ENV_CTRL_2,28,27);
  zz_decode_BRANCH_CTRL_1 <= zz_decode_BRANCH_CTRL_2;
  zz_decode_ENV_CTRL_9 <= pkg_extract(zz_decode_ENV_CTRL_2,30,30);
  zz_decode_ENV_CTRL_1 <= zz_decode_ENV_CTRL_9;
  decodeExceptionPort_valid <= (decode_arbitration_isValid and (not decode_LEGAL_INSTRUCTION));
  decodeExceptionPort_payload_code <= pkg_unsigned("0010");
  decodeExceptionPort_payload_badAddr <= unsigned(decode_INSTRUCTION);
  when_RegFilePlugin_l63 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,11,7) = pkg_stdLogicVector("00000"));
  decode_RegFilePlugin_regFileReadAddress1 <= unsigned(pkg_extract(decode_INSTRUCTION_ANTICIPATED,19,15));
  decode_RegFilePlugin_regFileReadAddress2 <= unsigned(pkg_extract(decode_INSTRUCTION_ANTICIPATED,24,20));
  decode_RegFilePlugin_rs1Data <= zz_RegFilePlugin_regFile_port0;
  decode_RegFilePlugin_rs2Data <= zz_RegFilePlugin_regFile_port0_1;
  process(zz_lastStageRegFileWrite_valid,writeBack_arbitration_isFiring,zz_3)
  begin
    lastStageRegFileWrite_valid <= (zz_lastStageRegFileWrite_valid and writeBack_arbitration_isFiring);
    if zz_3 = '1' then
      lastStageRegFileWrite_valid <= pkg_toStdLogic(true);
    end if;
  end process;

  process(zz_lastStageRegFileWrite_payload_address,zz_3)
  begin
    lastStageRegFileWrite_payload_address <= unsigned(pkg_extract(zz_lastStageRegFileWrite_payload_address,11,7));
    if zz_3 = '1' then
      lastStageRegFileWrite_payload_address <= pkg_unsigned("00000");
    end if;
  end process;

  process(zz_decode_RS2_2,zz_3)
  begin
    lastStageRegFileWrite_payload_data <= zz_decode_RS2_2;
    if zz_3 = '1' then
      lastStageRegFileWrite_payload_data <= pkg_stdLogicVector("00000000000000000000000000000000");
    end if;
  end process;

  process(execute_ALU_BITWISE_CTRL,execute_SRC1,execute_SRC2)
  begin
    case execute_ALU_BITWISE_CTRL is
      when AluBitwiseCtrlEnum_seq_AND_1 =>
        execute_IntAluPlugin_bitwise <= (execute_SRC1 and execute_SRC2);
      when AluBitwiseCtrlEnum_seq_OR_1 =>
        execute_IntAluPlugin_bitwise <= (execute_SRC1 or execute_SRC2);
      when others =>
        execute_IntAluPlugin_bitwise <= (execute_SRC1 xor execute_SRC2);
    end case;
  end process;

  process(execute_ALU_CTRL,execute_IntAluPlugin_bitwise,execute_SRC_LESS,execute_SRC_ADD_SUB)
  begin
    case execute_ALU_CTRL is
      when AluCtrlEnum_seq_BITWISE =>
        zz_execute_REGFILE_WRITE_DATA <= execute_IntAluPlugin_bitwise;
      when AluCtrlEnum_seq_SLT_SLTU =>
        zz_execute_REGFILE_WRITE_DATA <= pkg_resize(pkg_toStdLogicVector(execute_SRC_LESS),32);
      when others =>
        zz_execute_REGFILE_WRITE_DATA <= execute_SRC_ADD_SUB;
    end case;
  end process;

  process(execute_SRC1_CTRL,execute_RS1,execute_INSTRUCTION)
  begin
    case execute_SRC1_CTRL is
      when Src1CtrlEnum_seq_RS =>
        zz_execute_SRC1 <= execute_RS1;
      when Src1CtrlEnum_seq_PC_INCREMENT =>
        zz_execute_SRC1 <= pkg_resize(pkg_stdLogicVector("100"),32);
      when Src1CtrlEnum_seq_IMU =>
        zz_execute_SRC1 <= pkg_cat(pkg_extract(execute_INSTRUCTION,31,12),std_logic_vector(pkg_unsigned("000000000000")));
      when others =>
        zz_execute_SRC1 <= pkg_resize(pkg_extract(execute_INSTRUCTION,19,15),32);
    end case;
  end process;

  zz_execute_SRC2_1 <= pkg_extract(execute_INSTRUCTION,31);
  process(zz_execute_SRC2_1)
  begin
    zz_execute_SRC2_2(19) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(18) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(17) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(16) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(15) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(14) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(13) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(12) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(11) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(10) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(9) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(8) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(7) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(6) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(5) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(4) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(3) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(2) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(1) <= zz_execute_SRC2_1;
    zz_execute_SRC2_2(0) <= zz_execute_SRC2_1;
  end process;

  zz_execute_SRC2_3 <= pkg_extract(pkg_cat(pkg_extract(execute_INSTRUCTION,31,25),pkg_extract(execute_INSTRUCTION,11,7)),11);
  process(zz_execute_SRC2_3)
  begin
    zz_execute_SRC2_4(19) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(18) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(17) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(16) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(15) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(14) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(13) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(12) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(11) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(10) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(9) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(8) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(7) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(6) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(5) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(4) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(3) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(2) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(1) <= zz_execute_SRC2_3;
    zz_execute_SRC2_4(0) <= zz_execute_SRC2_3;
  end process;

  process(execute_SRC2_CTRL,execute_RS2,zz_execute_SRC2_2,execute_INSTRUCTION,zz_execute_SRC2_4,zz_execute_SRC2)
  begin
    case execute_SRC2_CTRL is
      when Src2CtrlEnum_seq_RS =>
        zz_execute_SRC2_5 <= execute_RS2;
      when Src2CtrlEnum_seq_IMI =>
        zz_execute_SRC2_5 <= pkg_cat(zz_execute_SRC2_2,pkg_extract(execute_INSTRUCTION,31,20));
      when Src2CtrlEnum_seq_IMS =>
        zz_execute_SRC2_5 <= pkg_cat(zz_execute_SRC2_4,pkg_cat(pkg_extract(execute_INSTRUCTION,31,25),pkg_extract(execute_INSTRUCTION,11,7)));
      when others =>
        zz_execute_SRC2_5 <= std_logic_vector(zz_execute_SRC2);
    end case;
  end process;

  process(execute_SRC1,execute_SRC_USE_SUB_LESS,execute_SRC2,execute_SRC2_FORCE_ZERO)
  begin
    execute_SrcPlugin_addSub <= std_logic_vector(((signed(execute_SRC1) + signed(pkg_mux(execute_SRC_USE_SUB_LESS,pkg_not(execute_SRC2),execute_SRC2))) + pkg_mux(execute_SRC_USE_SUB_LESS,pkg_signed("00000000000000000000000000000001"),pkg_signed("00000000000000000000000000000000"))));
    if execute_SRC2_FORCE_ZERO = '1' then
      execute_SrcPlugin_addSub <= execute_SRC1;
    end if;
  end process;

  execute_SrcPlugin_less <= pkg_mux(pkg_toStdLogic(pkg_extract(execute_SRC1,31) = pkg_extract(execute_SRC2,31)),pkg_extract(execute_SrcPlugin_addSub,31),pkg_mux(execute_SRC_LESS_UNSIGNED,pkg_extract(execute_SRC2,31),pkg_extract(execute_SRC1,31)));
  execute_FullBarrelShifterPlugin_amplitude <= unsigned(pkg_extract(execute_SRC2,4,0));
  process(execute_SRC1)
  begin
    zz_execute_FullBarrelShifterPlugin_reversed(0) <= pkg_extract(execute_SRC1,31);
    zz_execute_FullBarrelShifterPlugin_reversed(1) <= pkg_extract(execute_SRC1,30);
    zz_execute_FullBarrelShifterPlugin_reversed(2) <= pkg_extract(execute_SRC1,29);
    zz_execute_FullBarrelShifterPlugin_reversed(3) <= pkg_extract(execute_SRC1,28);
    zz_execute_FullBarrelShifterPlugin_reversed(4) <= pkg_extract(execute_SRC1,27);
    zz_execute_FullBarrelShifterPlugin_reversed(5) <= pkg_extract(execute_SRC1,26);
    zz_execute_FullBarrelShifterPlugin_reversed(6) <= pkg_extract(execute_SRC1,25);
    zz_execute_FullBarrelShifterPlugin_reversed(7) <= pkg_extract(execute_SRC1,24);
    zz_execute_FullBarrelShifterPlugin_reversed(8) <= pkg_extract(execute_SRC1,23);
    zz_execute_FullBarrelShifterPlugin_reversed(9) <= pkg_extract(execute_SRC1,22);
    zz_execute_FullBarrelShifterPlugin_reversed(10) <= pkg_extract(execute_SRC1,21);
    zz_execute_FullBarrelShifterPlugin_reversed(11) <= pkg_extract(execute_SRC1,20);
    zz_execute_FullBarrelShifterPlugin_reversed(12) <= pkg_extract(execute_SRC1,19);
    zz_execute_FullBarrelShifterPlugin_reversed(13) <= pkg_extract(execute_SRC1,18);
    zz_execute_FullBarrelShifterPlugin_reversed(14) <= pkg_extract(execute_SRC1,17);
    zz_execute_FullBarrelShifterPlugin_reversed(15) <= pkg_extract(execute_SRC1,16);
    zz_execute_FullBarrelShifterPlugin_reversed(16) <= pkg_extract(execute_SRC1,15);
    zz_execute_FullBarrelShifterPlugin_reversed(17) <= pkg_extract(execute_SRC1,14);
    zz_execute_FullBarrelShifterPlugin_reversed(18) <= pkg_extract(execute_SRC1,13);
    zz_execute_FullBarrelShifterPlugin_reversed(19) <= pkg_extract(execute_SRC1,12);
    zz_execute_FullBarrelShifterPlugin_reversed(20) <= pkg_extract(execute_SRC1,11);
    zz_execute_FullBarrelShifterPlugin_reversed(21) <= pkg_extract(execute_SRC1,10);
    zz_execute_FullBarrelShifterPlugin_reversed(22) <= pkg_extract(execute_SRC1,9);
    zz_execute_FullBarrelShifterPlugin_reversed(23) <= pkg_extract(execute_SRC1,8);
    zz_execute_FullBarrelShifterPlugin_reversed(24) <= pkg_extract(execute_SRC1,7);
    zz_execute_FullBarrelShifterPlugin_reversed(25) <= pkg_extract(execute_SRC1,6);
    zz_execute_FullBarrelShifterPlugin_reversed(26) <= pkg_extract(execute_SRC1,5);
    zz_execute_FullBarrelShifterPlugin_reversed(27) <= pkg_extract(execute_SRC1,4);
    zz_execute_FullBarrelShifterPlugin_reversed(28) <= pkg_extract(execute_SRC1,3);
    zz_execute_FullBarrelShifterPlugin_reversed(29) <= pkg_extract(execute_SRC1,2);
    zz_execute_FullBarrelShifterPlugin_reversed(30) <= pkg_extract(execute_SRC1,1);
    zz_execute_FullBarrelShifterPlugin_reversed(31) <= pkg_extract(execute_SRC1,0);
  end process;

  execute_FullBarrelShifterPlugin_reversed <= pkg_mux(pkg_toStdLogic(execute_SHIFT_CTRL = ShiftCtrlEnum_seq_SLL_1),zz_execute_FullBarrelShifterPlugin_reversed,execute_SRC1);
  process(execute_SHIFT_RIGHT)
  begin
    zz_decode_RS2_3(0) <= pkg_extract(execute_SHIFT_RIGHT,31);
    zz_decode_RS2_3(1) <= pkg_extract(execute_SHIFT_RIGHT,30);
    zz_decode_RS2_3(2) <= pkg_extract(execute_SHIFT_RIGHT,29);
    zz_decode_RS2_3(3) <= pkg_extract(execute_SHIFT_RIGHT,28);
    zz_decode_RS2_3(4) <= pkg_extract(execute_SHIFT_RIGHT,27);
    zz_decode_RS2_3(5) <= pkg_extract(execute_SHIFT_RIGHT,26);
    zz_decode_RS2_3(6) <= pkg_extract(execute_SHIFT_RIGHT,25);
    zz_decode_RS2_3(7) <= pkg_extract(execute_SHIFT_RIGHT,24);
    zz_decode_RS2_3(8) <= pkg_extract(execute_SHIFT_RIGHT,23);
    zz_decode_RS2_3(9) <= pkg_extract(execute_SHIFT_RIGHT,22);
    zz_decode_RS2_3(10) <= pkg_extract(execute_SHIFT_RIGHT,21);
    zz_decode_RS2_3(11) <= pkg_extract(execute_SHIFT_RIGHT,20);
    zz_decode_RS2_3(12) <= pkg_extract(execute_SHIFT_RIGHT,19);
    zz_decode_RS2_3(13) <= pkg_extract(execute_SHIFT_RIGHT,18);
    zz_decode_RS2_3(14) <= pkg_extract(execute_SHIFT_RIGHT,17);
    zz_decode_RS2_3(15) <= pkg_extract(execute_SHIFT_RIGHT,16);
    zz_decode_RS2_3(16) <= pkg_extract(execute_SHIFT_RIGHT,15);
    zz_decode_RS2_3(17) <= pkg_extract(execute_SHIFT_RIGHT,14);
    zz_decode_RS2_3(18) <= pkg_extract(execute_SHIFT_RIGHT,13);
    zz_decode_RS2_3(19) <= pkg_extract(execute_SHIFT_RIGHT,12);
    zz_decode_RS2_3(20) <= pkg_extract(execute_SHIFT_RIGHT,11);
    zz_decode_RS2_3(21) <= pkg_extract(execute_SHIFT_RIGHT,10);
    zz_decode_RS2_3(22) <= pkg_extract(execute_SHIFT_RIGHT,9);
    zz_decode_RS2_3(23) <= pkg_extract(execute_SHIFT_RIGHT,8);
    zz_decode_RS2_3(24) <= pkg_extract(execute_SHIFT_RIGHT,7);
    zz_decode_RS2_3(25) <= pkg_extract(execute_SHIFT_RIGHT,6);
    zz_decode_RS2_3(26) <= pkg_extract(execute_SHIFT_RIGHT,5);
    zz_decode_RS2_3(27) <= pkg_extract(execute_SHIFT_RIGHT,4);
    zz_decode_RS2_3(28) <= pkg_extract(execute_SHIFT_RIGHT,3);
    zz_decode_RS2_3(29) <= pkg_extract(execute_SHIFT_RIGHT,2);
    zz_decode_RS2_3(30) <= pkg_extract(execute_SHIFT_RIGHT,1);
    zz_decode_RS2_3(31) <= pkg_extract(execute_SHIFT_RIGHT,0);
  end process;

  execute_MulPlugin_a <= execute_RS1;
  execute_MulPlugin_b <= execute_RS2;
  switch_MulPlugin_l87 <= pkg_extract(execute_INSTRUCTION,13,12);
  process(switch_MulPlugin_l87)
  begin
    case switch_MulPlugin_l87 is
      when "01" =>
        execute_MulPlugin_aSigned <= pkg_toStdLogic(true);
      when "10" =>
        execute_MulPlugin_aSigned <= pkg_toStdLogic(true);
      when others =>
        execute_MulPlugin_aSigned <= pkg_toStdLogic(false);
    end case;
  end process;

  process(switch_MulPlugin_l87)
  begin
    case switch_MulPlugin_l87 is
      when "01" =>
        execute_MulPlugin_bSigned <= pkg_toStdLogic(true);
      when "10" =>
        execute_MulPlugin_bSigned <= pkg_toStdLogic(false);
      when others =>
        execute_MulPlugin_bSigned <= pkg_toStdLogic(false);
    end case;
  end process;

  execute_MulPlugin_aULow <= unsigned(pkg_extract(execute_MulPlugin_a,15,0));
  execute_MulPlugin_bULow <= unsigned(pkg_extract(execute_MulPlugin_b,15,0));
  execute_MulPlugin_aSLow <= signed(pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(false)),pkg_extract(execute_MulPlugin_a,15,0)));
  execute_MulPlugin_bSLow <= signed(pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic(false)),pkg_extract(execute_MulPlugin_b,15,0)));
  execute_MulPlugin_aHigh <= signed(pkg_cat(pkg_toStdLogicVector((execute_MulPlugin_aSigned and pkg_extract(execute_MulPlugin_a,31))),pkg_extract(execute_MulPlugin_a,31,16)));
  execute_MulPlugin_bHigh <= signed(pkg_cat(pkg_toStdLogicVector((execute_MulPlugin_bSigned and pkg_extract(execute_MulPlugin_b,31))),pkg_extract(execute_MulPlugin_b,31,16)));
  writeBack_MulPlugin_result <= (pkg_resize(writeBack_MUL_LOW,66) + pkg_shiftLeft(writeBack_MUL_HH,32));
  when_MulPlugin_l147 <= (writeBack_arbitration_isValid and writeBack_IS_MUL);
  switch_MulPlugin_l148 <= pkg_extract(writeBack_INSTRUCTION,13,12);
  memory_DivPlugin_frontendOk <= pkg_toStdLogic(true);
  process(when_MulDivIterativePlugin_l128,when_MulDivIterativePlugin_l132)
  begin
    memory_DivPlugin_div_counter_willIncrement <= pkg_toStdLogic(false);
    if when_MulDivIterativePlugin_l128 = '1' then
      if when_MulDivIterativePlugin_l132 = '1' then
        memory_DivPlugin_div_counter_willIncrement <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  process(when_MulDivIterativePlugin_l162)
  begin
    memory_DivPlugin_div_counter_willClear <= pkg_toStdLogic(false);
    if when_MulDivIterativePlugin_l162 = '1' then
      memory_DivPlugin_div_counter_willClear <= pkg_toStdLogic(true);
    end if;
  end process;

  memory_DivPlugin_div_counter_willOverflowIfInc <= pkg_toStdLogic(memory_DivPlugin_div_counter_value = pkg_unsigned("100001"));
  memory_DivPlugin_div_counter_willOverflow <= (memory_DivPlugin_div_counter_willOverflowIfInc and memory_DivPlugin_div_counter_willIncrement);
  process(memory_DivPlugin_div_counter_willOverflow,memory_DivPlugin_div_counter_value,memory_DivPlugin_div_counter_willIncrement,memory_DivPlugin_div_counter_willClear)
  begin
    if memory_DivPlugin_div_counter_willOverflow = '1' then
      memory_DivPlugin_div_counter_valueNext <= pkg_unsigned("000000");
    else
      memory_DivPlugin_div_counter_valueNext <= (memory_DivPlugin_div_counter_value + pkg_resize(unsigned(pkg_toStdLogicVector(memory_DivPlugin_div_counter_willIncrement)),6));
    end if;
    if memory_DivPlugin_div_counter_willClear = '1' then
      memory_DivPlugin_div_counter_valueNext <= pkg_unsigned("000000");
    end if;
  end process;

  when_MulDivIterativePlugin_l126 <= pkg_toStdLogic(memory_DivPlugin_div_counter_value = pkg_unsigned("100000"));
  when_MulDivIterativePlugin_l126_1 <= (not memory_arbitration_isStuck);
  when_MulDivIterativePlugin_l128 <= (memory_arbitration_isValid and memory_IS_DIV);
  when_MulDivIterativePlugin_l129 <= ((not memory_DivPlugin_frontendOk) or (not memory_DivPlugin_div_done));
  when_MulDivIterativePlugin_l132 <= (memory_DivPlugin_frontendOk and (not memory_DivPlugin_div_done));
  zz_memory_DivPlugin_div_stage_0_remainderShifted <= pkg_extract(memory_DivPlugin_rs1,31,0);
  memory_DivPlugin_div_stage_0_remainderShifted <= unsigned(pkg_cat(std_logic_vector(pkg_extract(memory_DivPlugin_accumulator,31,0)),pkg_toStdLogicVector(pkg_extract(zz_memory_DivPlugin_div_stage_0_remainderShifted,31))));
  memory_DivPlugin_div_stage_0_remainderMinusDenominator <= (memory_DivPlugin_div_stage_0_remainderShifted - pkg_resize(memory_DivPlugin_rs2,33));
  memory_DivPlugin_div_stage_0_outRemainder <= pkg_mux((not pkg_extract(memory_DivPlugin_div_stage_0_remainderMinusDenominator,32)),pkg_resize(memory_DivPlugin_div_stage_0_remainderMinusDenominator,32),pkg_resize(memory_DivPlugin_div_stage_0_remainderShifted,32));
  memory_DivPlugin_div_stage_0_outNumerator <= pkg_resize(unsigned(pkg_cat(std_logic_vector(zz_memory_DivPlugin_div_stage_0_remainderShifted),pkg_toStdLogicVector((not pkg_extract(memory_DivPlugin_div_stage_0_remainderMinusDenominator,32))))),32);
  when_MulDivIterativePlugin_l151 <= pkg_toStdLogic(memory_DivPlugin_div_counter_value = pkg_unsigned("100000"));
  zz_memory_DivPlugin_div_result <= pkg_mux(pkg_extract(memory_INSTRUCTION,13),pkg_extract(memory_DivPlugin_accumulator,31,0),pkg_extract(memory_DivPlugin_rs1,31,0));
  when_MulDivIterativePlugin_l162 <= (not memory_arbitration_isStuck);
  zz_memory_DivPlugin_rs2 <= (pkg_extract(execute_RS2,31) and execute_IS_RS2_SIGNED);
  zz_memory_DivPlugin_rs1 <= (pkg_toStdLogic(false) or ((execute_IS_DIV and pkg_extract(execute_RS1,31)) and execute_IS_RS1_SIGNED));
  process(execute_IS_RS1_SIGNED,execute_RS1)
  begin
    zz_memory_DivPlugin_rs1_1(32) <= (execute_IS_RS1_SIGNED and pkg_extract(execute_RS1,31));
    zz_memory_DivPlugin_rs1_1(31 downto 0) <= execute_RS1;
  end process;

  process(when_HazardSimplePlugin_l57,when_HazardSimplePlugin_l58,when_HazardSimplePlugin_l48,when_HazardSimplePlugin_l57_1,when_HazardSimplePlugin_l58_1,when_HazardSimplePlugin_l48_1,when_HazardSimplePlugin_l57_2,when_HazardSimplePlugin_l58_2,when_HazardSimplePlugin_l48_2,when_HazardSimplePlugin_l105)
  begin
    HazardSimplePlugin_src0Hazard <= pkg_toStdLogic(false);
    if when_HazardSimplePlugin_l57 = '1' then
      if when_HazardSimplePlugin_l58 = '1' then
        if when_HazardSimplePlugin_l48 = '1' then
          HazardSimplePlugin_src0Hazard <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l57_1 = '1' then
      if when_HazardSimplePlugin_l58_1 = '1' then
        if when_HazardSimplePlugin_l48_1 = '1' then
          HazardSimplePlugin_src0Hazard <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l57_2 = '1' then
      if when_HazardSimplePlugin_l58_2 = '1' then
        if when_HazardSimplePlugin_l48_2 = '1' then
          HazardSimplePlugin_src0Hazard <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l105 = '1' then
      HazardSimplePlugin_src0Hazard <= pkg_toStdLogic(false);
    end if;
  end process;

  process(when_HazardSimplePlugin_l57,when_HazardSimplePlugin_l58,when_HazardSimplePlugin_l51,when_HazardSimplePlugin_l57_1,when_HazardSimplePlugin_l58_1,when_HazardSimplePlugin_l51_1,when_HazardSimplePlugin_l57_2,when_HazardSimplePlugin_l58_2,when_HazardSimplePlugin_l51_2,when_HazardSimplePlugin_l108)
  begin
    HazardSimplePlugin_src1Hazard <= pkg_toStdLogic(false);
    if when_HazardSimplePlugin_l57 = '1' then
      if when_HazardSimplePlugin_l58 = '1' then
        if when_HazardSimplePlugin_l51 = '1' then
          HazardSimplePlugin_src1Hazard <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l57_1 = '1' then
      if when_HazardSimplePlugin_l58_1 = '1' then
        if when_HazardSimplePlugin_l51_1 = '1' then
          HazardSimplePlugin_src1Hazard <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l57_2 = '1' then
      if when_HazardSimplePlugin_l58_2 = '1' then
        if when_HazardSimplePlugin_l51_2 = '1' then
          HazardSimplePlugin_src1Hazard <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
    if when_HazardSimplePlugin_l108 = '1' then
      HazardSimplePlugin_src1Hazard <= pkg_toStdLogic(false);
    end if;
  end process;

  HazardSimplePlugin_writeBackWrites_valid <= (zz_lastStageRegFileWrite_valid and writeBack_arbitration_isFiring);
  HazardSimplePlugin_writeBackWrites_payload_address <= pkg_extract(zz_lastStageRegFileWrite_payload_address,11,7);
  HazardSimplePlugin_writeBackWrites_payload_data <= zz_decode_RS2_2;
  HazardSimplePlugin_addr0Match <= pkg_toStdLogic(HazardSimplePlugin_writeBackBuffer_payload_address = pkg_extract(decode_INSTRUCTION,19,15));
  HazardSimplePlugin_addr1Match <= pkg_toStdLogic(HazardSimplePlugin_writeBackBuffer_payload_address = pkg_extract(decode_INSTRUCTION,24,20));
  when_HazardSimplePlugin_l47 <= pkg_toStdLogic(true);
  when_HazardSimplePlugin_l48 <= pkg_toStdLogic(pkg_extract(writeBack_INSTRUCTION,11,7) = pkg_extract(decode_INSTRUCTION,19,15));
  when_HazardSimplePlugin_l51 <= pkg_toStdLogic(pkg_extract(writeBack_INSTRUCTION,11,7) = pkg_extract(decode_INSTRUCTION,24,20));
  when_HazardSimplePlugin_l45 <= (writeBack_arbitration_isValid and writeBack_REGFILE_WRITE_VALID);
  when_HazardSimplePlugin_l57 <= (writeBack_arbitration_isValid and writeBack_REGFILE_WRITE_VALID);
  when_HazardSimplePlugin_l58 <= (pkg_toStdLogic(false) or (not when_HazardSimplePlugin_l47));
  when_HazardSimplePlugin_l48_1 <= pkg_toStdLogic(pkg_extract(memory_INSTRUCTION,11,7) = pkg_extract(decode_INSTRUCTION,19,15));
  when_HazardSimplePlugin_l51_1 <= pkg_toStdLogic(pkg_extract(memory_INSTRUCTION,11,7) = pkg_extract(decode_INSTRUCTION,24,20));
  when_HazardSimplePlugin_l45_1 <= (memory_arbitration_isValid and memory_REGFILE_WRITE_VALID);
  when_HazardSimplePlugin_l57_1 <= (memory_arbitration_isValid and memory_REGFILE_WRITE_VALID);
  when_HazardSimplePlugin_l58_1 <= (pkg_toStdLogic(false) or (not memory_BYPASSABLE_MEMORY_STAGE));
  when_HazardSimplePlugin_l48_2 <= pkg_toStdLogic(pkg_extract(execute_INSTRUCTION,11,7) = pkg_extract(decode_INSTRUCTION,19,15));
  when_HazardSimplePlugin_l51_2 <= pkg_toStdLogic(pkg_extract(execute_INSTRUCTION,11,7) = pkg_extract(decode_INSTRUCTION,24,20));
  when_HazardSimplePlugin_l45_2 <= (execute_arbitration_isValid and execute_REGFILE_WRITE_VALID);
  when_HazardSimplePlugin_l57_2 <= (execute_arbitration_isValid and execute_REGFILE_WRITE_VALID);
  when_HazardSimplePlugin_l58_2 <= (pkg_toStdLogic(false) or (not execute_BYPASSABLE_EXECUTE_STAGE));
  when_HazardSimplePlugin_l105 <= (not decode_RS1_USE);
  when_HazardSimplePlugin_l108 <= (not decode_RS2_USE);
  when_HazardSimplePlugin_l113 <= (decode_arbitration_isValid and (HazardSimplePlugin_src0Hazard or HazardSimplePlugin_src1Hazard));
  execute_BranchPlugin_eq <= pkg_toStdLogic(execute_SRC1 = execute_SRC2);
  switch_Misc_l204_1 <= pkg_extract(execute_INSTRUCTION,14,12);
  process(switch_Misc_l204_1,execute_BranchPlugin_eq,execute_SRC_LESS)
  begin
    if (switch_Misc_l204_1 = pkg_stdLogicVector("000")) then
        zz_execute_BRANCH_DO <= execute_BranchPlugin_eq;
    elsif (switch_Misc_l204_1 = pkg_stdLogicVector("001")) then
        zz_execute_BRANCH_DO <= (not execute_BranchPlugin_eq);
    elsif (pkg_toStdLogic((switch_Misc_l204_1 and pkg_stdLogicVector("101")) = pkg_stdLogicVector("101")) = '1') then
        zz_execute_BRANCH_DO <= (not execute_SRC_LESS);
    else
        zz_execute_BRANCH_DO <= execute_SRC_LESS;
    end if;
  end process;

  process(execute_BRANCH_CTRL,zz_execute_BRANCH_DO)
  begin
    case execute_BRANCH_CTRL is
      when BranchCtrlEnum_seq_INC =>
        zz_execute_BRANCH_DO_1 <= pkg_toStdLogic(false);
      when BranchCtrlEnum_seq_JAL =>
        zz_execute_BRANCH_DO_1 <= pkg_toStdLogic(true);
      when BranchCtrlEnum_seq_JALR =>
        zz_execute_BRANCH_DO_1 <= pkg_toStdLogic(true);
      when others =>
        zz_execute_BRANCH_DO_1 <= zz_execute_BRANCH_DO;
    end case;
  end process;

  execute_BranchPlugin_branch_src1 <= pkg_mux(pkg_toStdLogic(execute_BRANCH_CTRL = BranchCtrlEnum_seq_JALR),unsigned(execute_RS1),execute_PC);
  zz_execute_BRANCH_SRC22 <= pkg_extract(pkg_cat(pkg_cat(pkg_cat(pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,31)),pkg_extract(execute_INSTRUCTION,19,12)),pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,20))),pkg_extract(execute_INSTRUCTION,30,21)),19);
  process(zz_execute_BRANCH_SRC22)
  begin
    zz_execute_BRANCH_SRC22_1(10) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(9) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(8) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(7) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(6) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(5) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(4) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(3) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(2) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(1) <= zz_execute_BRANCH_SRC22;
    zz_execute_BRANCH_SRC22_1(0) <= zz_execute_BRANCH_SRC22;
  end process;

  zz_execute_BRANCH_SRC22_2 <= pkg_extract(execute_INSTRUCTION,31);
  process(zz_execute_BRANCH_SRC22_2)
  begin
    zz_execute_BRANCH_SRC22_3(19) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(18) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(17) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(16) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(15) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(14) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(13) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(12) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(11) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(10) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(9) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(8) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(7) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(6) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(5) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(4) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(3) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(2) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(1) <= zz_execute_BRANCH_SRC22_2;
    zz_execute_BRANCH_SRC22_3(0) <= zz_execute_BRANCH_SRC22_2;
  end process;

  zz_execute_BRANCH_SRC22_4 <= pkg_extract(pkg_cat(pkg_cat(pkg_cat(pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,31)),pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,7))),pkg_extract(execute_INSTRUCTION,30,25)),pkg_extract(execute_INSTRUCTION,11,8)),11);
  process(zz_execute_BRANCH_SRC22_4)
  begin
    zz_execute_BRANCH_SRC22_5(18) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(17) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(16) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(15) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(14) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(13) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(12) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(11) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(10) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(9) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(8) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(7) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(6) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(5) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(4) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(3) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(2) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(1) <= zz_execute_BRANCH_SRC22_4;
    zz_execute_BRANCH_SRC22_5(0) <= zz_execute_BRANCH_SRC22_4;
  end process;

  process(execute_BRANCH_CTRL,zz_execute_BRANCH_SRC22_1,execute_INSTRUCTION,zz_execute_BRANCH_SRC22_3,zz_execute_BRANCH_SRC22_5)
  begin
    case execute_BRANCH_CTRL is
      when BranchCtrlEnum_seq_JAL =>
        zz_execute_BRANCH_SRC22_6 <= pkg_cat(pkg_cat(zz_execute_BRANCH_SRC22_1,pkg_cat(pkg_cat(pkg_cat(pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,31)),pkg_extract(execute_INSTRUCTION,19,12)),pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,20))),pkg_extract(execute_INSTRUCTION,30,21))),pkg_toStdLogicVector(pkg_toStdLogic(false)));
      when BranchCtrlEnum_seq_JALR =>
        zz_execute_BRANCH_SRC22_6 <= pkg_cat(zz_execute_BRANCH_SRC22_3,pkg_extract(execute_INSTRUCTION,31,20));
      when others =>
        zz_execute_BRANCH_SRC22_6 <= pkg_cat(pkg_cat(zz_execute_BRANCH_SRC22_5,pkg_cat(pkg_cat(pkg_cat(pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,31)),pkg_toStdLogicVector(pkg_extract(execute_INSTRUCTION,7))),pkg_extract(execute_INSTRUCTION,30,25)),pkg_extract(execute_INSTRUCTION,11,8))),pkg_toStdLogicVector(pkg_toStdLogic(false)));
    end case;
  end process;

  execute_BranchPlugin_branchAdder <= (execute_BranchPlugin_branch_src1 + execute_BRANCH_SRC22);
  memory_BranchPlugin_predictionMissmatch <= (pkg_toStdLogic(IBusCachedPlugin_fetchPrediction_cmd_hadBranch /= memory_BRANCH_DO) or (memory_BRANCH_DO and memory_TARGET_MISSMATCH2));
  IBusCachedPlugin_fetchPrediction_rsp_wasRight <= (not memory_BranchPlugin_predictionMissmatch);
  IBusCachedPlugin_fetchPrediction_rsp_finalPc <= memory_BRANCH_CALC;
  IBusCachedPlugin_fetchPrediction_rsp_sourceLastWord <= memory_PC;
  BranchPlugin_jumpInterface_valid <= ((memory_arbitration_isValid and memory_BranchPlugin_predictionMissmatch) and (not pkg_toStdLogic(false)));
  BranchPlugin_jumpInterface_payload <= pkg_mux(memory_BRANCH_DO,memory_BRANCH_CALC,memory_NEXT_PC2);
  BranchPlugin_branchExceptionPort_valid <= ((memory_arbitration_isValid and memory_BRANCH_DO) and pkg_extract(memory_BRANCH_CALC,1));
  BranchPlugin_branchExceptionPort_payload_code <= pkg_unsigned("0000");
  BranchPlugin_branchExceptionPort_payload_badAddr <= memory_BRANCH_CALC;
  process(CsrPlugin_forceMachineWire)
  begin
    CsrPlugin_privilege <= pkg_unsigned("11");
    if CsrPlugin_forceMachineWire = '1' then
      CsrPlugin_privilege <= pkg_unsigned("11");
    end if;
  end process;

  CsrPlugin_misa_base <= pkg_unsigned("01");
  CsrPlugin_misa_extensions <= pkg_stdLogicVector("00000000000000000001000010");
  CsrPlugin_mtvec_mode <= pkg_stdLogicVector("00");
  CsrPlugin_mtvec_base <= pkg_unsigned("000000000000000000000000001000");
  zz_when_CsrPlugin_l952 <= (CsrPlugin_mip_MTIP and CsrPlugin_mie_MTIE);
  zz_when_CsrPlugin_l952_1 <= (CsrPlugin_mip_MSIP and CsrPlugin_mie_MSIE);
  zz_when_CsrPlugin_l952_2 <= (CsrPlugin_mip_MEIP and CsrPlugin_mie_MEIE);
  CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped <= pkg_unsigned("11");
  CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege <= pkg_mux(pkg_toStdLogic(CsrPlugin_privilege < CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped),CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped,CsrPlugin_privilege);
  zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code <= unsigned(pkg_cat(pkg_toStdLogicVector(decodeExceptionPort_valid),pkg_toStdLogicVector(IBusCachedPlugin_decodeExceptionPort_valid)));
  zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 <= pkg_extract(std_logic_vector((zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code and pkg_not((zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code - pkg_unsigned("01"))))),0);
  process(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode,zz_when,decode_arbitration_isFlushed)
  begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_decode <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
    if zz_when = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode <= pkg_toStdLogic(true);
    end if;
    if decode_arbitration_isFlushed = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode <= pkg_toStdLogic(false);
    end if;
  end process;

  process(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute,execute_arbitration_isFlushed)
  begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_execute <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
    if execute_arbitration_isFlushed = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute <= pkg_toStdLogic(false);
    end if;
  end process;

  process(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory,BranchPlugin_branchExceptionPort_valid,memory_arbitration_isFlushed)
  begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_memory <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
    if BranchPlugin_branchExceptionPort_valid = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory <= pkg_toStdLogic(true);
    end if;
    if memory_arbitration_isFlushed = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory <= pkg_toStdLogic(false);
    end if;
  end process;

  process(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack,DBusCachedPlugin_exceptionBus_valid,writeBack_arbitration_isFlushed)
  begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
    if DBusCachedPlugin_exceptionBus_valid = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack <= pkg_toStdLogic(true);
    end if;
    if writeBack_arbitration_isFlushed = '1' then
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack <= pkg_toStdLogic(false);
    end if;
  end process;

  when_CsrPlugin_l909 <= (not decode_arbitration_isStuck);
  when_CsrPlugin_l909_1 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l909_2 <= (not memory_arbitration_isStuck);
  when_CsrPlugin_l909_3 <= (not writeBack_arbitration_isStuck);
  when_CsrPlugin_l922 <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack),pkg_cat(pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValids_memory),pkg_cat(pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValids_execute),pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValids_decode)))) /= pkg_stdLogicVector("0000"));
  CsrPlugin_exceptionPendings_0 <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  CsrPlugin_exceptionPendings_1 <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  CsrPlugin_exceptionPendings_2 <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  CsrPlugin_exceptionPendings_3 <= CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  when_CsrPlugin_l946 <= (CsrPlugin_mstatus_MIE or pkg_toStdLogic(CsrPlugin_privilege < pkg_unsigned("11")));
  when_CsrPlugin_l952 <= ((zz_when_CsrPlugin_l952 and pkg_toStdLogic(true)) and (not pkg_toStdLogic(false)));
  when_CsrPlugin_l952_1 <= ((zz_when_CsrPlugin_l952_1 and pkg_toStdLogic(true)) and (not pkg_toStdLogic(false)));
  when_CsrPlugin_l952_2 <= ((zz_when_CsrPlugin_l952_2 and pkg_toStdLogic(true)) and (not pkg_toStdLogic(false)));
  CsrPlugin_exception <= (CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack and CsrPlugin_allowException);
  CsrPlugin_lastStageWasWfi <= pkg_toStdLogic(false);
  CsrPlugin_pipelineLiberator_active <= ((CsrPlugin_interrupt_valid and CsrPlugin_allowInterrupts) and decode_arbitration_isValid);
  when_CsrPlugin_l980 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l980_1 <= (not memory_arbitration_isStuck);
  when_CsrPlugin_l980_2 <= (not writeBack_arbitration_isStuck);
  when_CsrPlugin_l985 <= ((not CsrPlugin_pipelineLiberator_active) or decode_arbitration_removeIt);
  process(CsrPlugin_pipelineLiberator_pcValids_2,when_CsrPlugin_l991,CsrPlugin_hadException)
  begin
    CsrPlugin_pipelineLiberator_done <= CsrPlugin_pipelineLiberator_pcValids_2;
    if when_CsrPlugin_l991 = '1' then
      CsrPlugin_pipelineLiberator_done <= pkg_toStdLogic(false);
    end if;
    if CsrPlugin_hadException = '1' then
      CsrPlugin_pipelineLiberator_done <= pkg_toStdLogic(false);
    end if;
  end process;

  when_CsrPlugin_l991 <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack),pkg_cat(pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory),pkg_toStdLogicVector(CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute))) /= pkg_stdLogicVector("000"));
  CsrPlugin_interruptJump <= ((CsrPlugin_interrupt_valid and CsrPlugin_pipelineLiberator_done) and CsrPlugin_allowInterrupts);
  process(CsrPlugin_interrupt_targetPrivilege,CsrPlugin_hadException,CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege)
  begin
    CsrPlugin_targetPrivilege <= CsrPlugin_interrupt_targetPrivilege;
    if CsrPlugin_hadException = '1' then
      CsrPlugin_targetPrivilege <= CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
    end if;
  end process;

  process(CsrPlugin_interrupt_code,CsrPlugin_hadException,CsrPlugin_exceptionPortCtrl_exceptionContext_code)
  begin
    CsrPlugin_trapCause <= pkg_resize(CsrPlugin_interrupt_code,4);
    if CsrPlugin_hadException = '1' then
      CsrPlugin_trapCause <= CsrPlugin_exceptionPortCtrl_exceptionContext_code;
    end if;
  end process;

  process(CsrPlugin_targetPrivilege,CsrPlugin_mtvec_mode)
  begin
    CsrPlugin_xtvec_mode <= pkg_stdLogicVector("XX");
    case CsrPlugin_targetPrivilege is
      when "11" =>
        CsrPlugin_xtvec_mode <= CsrPlugin_mtvec_mode;
      when others =>
    end case;
  end process;

  process(CsrPlugin_targetPrivilege,CsrPlugin_mtvec_base)
  begin
    CsrPlugin_xtvec_base <= pkg_unsigned("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
    case CsrPlugin_targetPrivilege is
      when "11" =>
        CsrPlugin_xtvec_base <= CsrPlugin_mtvec_base;
      when others =>
    end case;
  end process;

  when_CsrPlugin_l1019 <= (CsrPlugin_hadException or CsrPlugin_interruptJump);
  when_CsrPlugin_l1064 <= (writeBack_arbitration_isValid and pkg_toStdLogic(writeBack_ENV_CTRL = EnvCtrlEnum_seq_XRET));
  switch_CsrPlugin_l1068 <= pkg_extract(writeBack_INSTRUCTION,29,28);
  contextSwitching <= CsrPlugin_jumpInterface_valid;
  when_CsrPlugin_l1116 <= pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector((writeBack_arbitration_isValid and pkg_toStdLogic(writeBack_ENV_CTRL = EnvCtrlEnum_seq_XRET))),pkg_cat(pkg_toStdLogicVector((memory_arbitration_isValid and pkg_toStdLogic(memory_ENV_CTRL = EnvCtrlEnum_seq_XRET))),pkg_toStdLogicVector((execute_arbitration_isValid and pkg_toStdLogic(execute_ENV_CTRL = EnvCtrlEnum_seq_XRET))))) /= pkg_stdLogicVector("000"));
  execute_CsrPlugin_blockedBySideEffects <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_isValid),pkg_toStdLogicVector(memory_arbitration_isValid)) /= pkg_stdLogicVector("00")) or pkg_toStdLogic(false));
  process(execute_CsrPlugin_csr_768,execute_CsrPlugin_csr_836,execute_CsrPlugin_csr_772,execute_CsrPlugin_csr_833,execute_CsrPlugin_csr_834,execute_CSR_READ_OPCODE,execute_CsrPlugin_csr_835,CsrPlugin_csrMapping_allowCsrSignal,when_CsrPlugin_l1297,when_CsrPlugin_l1302)
  begin
    execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(true);
    if execute_CsrPlugin_csr_768 = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
    end if;
    if execute_CsrPlugin_csr_836 = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
    end if;
    if execute_CsrPlugin_csr_772 = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
    end if;
    if execute_CsrPlugin_csr_833 = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
    end if;
    if execute_CsrPlugin_csr_834 = '1' then
      if execute_CSR_READ_OPCODE = '1' then
        execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
      end if;
    end if;
    if execute_CsrPlugin_csr_835 = '1' then
      if execute_CSR_READ_OPCODE = '1' then
        execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
      end if;
    end if;
    if CsrPlugin_csrMapping_allowCsrSignal = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
    end if;
    if when_CsrPlugin_l1297 = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(true);
    end if;
    if when_CsrPlugin_l1302 = '1' then
      execute_CsrPlugin_illegalAccess <= pkg_toStdLogic(false);
    end if;
  end process;

  process(when_CsrPlugin_l1136,when_CsrPlugin_l1137)
  begin
    execute_CsrPlugin_illegalInstruction <= pkg_toStdLogic(false);
    if when_CsrPlugin_l1136 = '1' then
      if when_CsrPlugin_l1137 = '1' then
        execute_CsrPlugin_illegalInstruction <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  when_CsrPlugin_l1136 <= (execute_arbitration_isValid and pkg_toStdLogic(execute_ENV_CTRL = EnvCtrlEnum_seq_XRET));
  when_CsrPlugin_l1137 <= pkg_toStdLogic(CsrPlugin_privilege < unsigned(pkg_extract(execute_INSTRUCTION,29,28)));
  process(execute_arbitration_isValid,execute_IS_CSR,execute_CSR_WRITE_OPCODE,when_CsrPlugin_l1297)
  begin
    execute_CsrPlugin_writeInstruction <= ((execute_arbitration_isValid and execute_IS_CSR) and execute_CSR_WRITE_OPCODE);
    if when_CsrPlugin_l1297 = '1' then
      execute_CsrPlugin_writeInstruction <= pkg_toStdLogic(false);
    end if;
  end process;

  process(execute_arbitration_isValid,execute_IS_CSR,execute_CSR_READ_OPCODE,when_CsrPlugin_l1297)
  begin
    execute_CsrPlugin_readInstruction <= ((execute_arbitration_isValid and execute_IS_CSR) and execute_CSR_READ_OPCODE);
    if when_CsrPlugin_l1297 = '1' then
      execute_CsrPlugin_readInstruction <= pkg_toStdLogic(false);
    end if;
  end process;

  execute_CsrPlugin_writeEnable <= (execute_CsrPlugin_writeInstruction and (not execute_arbitration_isStuck));
  execute_CsrPlugin_readEnable <= (execute_CsrPlugin_readInstruction and (not execute_arbitration_isStuck));
  CsrPlugin_csrMapping_hazardFree <= (not execute_CsrPlugin_blockedBySideEffects);
  execute_CsrPlugin_readToWriteData <= CsrPlugin_csrMapping_readDataSignal;
  switch_Misc_l204_2 <= pkg_extract(execute_INSTRUCTION,13);
  process(switch_Misc_l204_2,execute_SRC1,execute_INSTRUCTION,execute_CsrPlugin_readToWriteData)
  begin
    case switch_Misc_l204_2 is
      when '0' =>
        zz_CsrPlugin_csrMapping_writeDataSignal <= execute_SRC1;
      when others =>
        zz_CsrPlugin_csrMapping_writeDataSignal <= pkg_mux(pkg_extract(execute_INSTRUCTION,12),(execute_CsrPlugin_readToWriteData and pkg_not(execute_SRC1)),(execute_CsrPlugin_readToWriteData or execute_SRC1));
    end case;
  end process;

  CsrPlugin_csrMapping_writeDataSignal <= zz_CsrPlugin_csrMapping_writeDataSignal;
  when_CsrPlugin_l1176 <= (execute_arbitration_isValid and execute_IS_CSR);
  when_CsrPlugin_l1180 <= (execute_arbitration_isValid and (execute_IS_CSR or pkg_toStdLogic(false)));
  execute_CsrPlugin_csrAddress <= pkg_extract(execute_INSTRUCTION,31,20);
  when_DebugPlugin_l225 <= (DebugPlugin_haltIt and (not DebugPlugin_isPipBusy));
  DebugPlugin_allowEBreak <= (DebugPlugin_debugUsed and (not DebugPlugin_disableEbreak));
  process(debug_bus_cmd_valid,switch_DebugPlugin_l267,debug_bus_cmd_payload_wr,IBusCachedPlugin_injectionPort_ready)
  begin
    debug_bus_cmd_ready_read_buffer <= pkg_toStdLogic(true);
    if debug_bus_cmd_valid = '1' then
      case switch_DebugPlugin_l267 is
        when "000001" =>
          if debug_bus_cmd_payload_wr = '1' then
            debug_bus_cmd_ready_read_buffer <= IBusCachedPlugin_injectionPort_ready;
          end if;
        when others =>
      end case;
    end if;
  end process;

  process(DebugPlugin_busReadDataReg,when_DebugPlugin_l244,DebugPlugin_resetIt,DebugPlugin_haltIt,DebugPlugin_isPipBusy,DebugPlugin_haltedByBreak,DebugPlugin_stepIt)
  begin
    debug_bus_rsp_data <= DebugPlugin_busReadDataReg;
    if when_DebugPlugin_l244 = '1' then
      debug_bus_rsp_data(0) <= DebugPlugin_resetIt;
      debug_bus_rsp_data(1) <= DebugPlugin_haltIt;
      debug_bus_rsp_data(2) <= DebugPlugin_isPipBusy;
      debug_bus_rsp_data(3) <= DebugPlugin_haltedByBreak;
      debug_bus_rsp_data(4) <= DebugPlugin_stepIt;
    end if;
  end process;

  when_DebugPlugin_l244 <= (not zz_when_DebugPlugin_l244);
  process(debug_bus_cmd_valid,switch_DebugPlugin_l267,debug_bus_cmd_payload_wr)
  begin
    IBusCachedPlugin_injectionPort_valid <= pkg_toStdLogic(false);
    if debug_bus_cmd_valid = '1' then
      case switch_DebugPlugin_l267 is
        when "000001" =>
          if debug_bus_cmd_payload_wr = '1' then
            IBusCachedPlugin_injectionPort_valid <= pkg_toStdLogic(true);
          end if;
        when others =>
      end case;
    end if;
  end process;

  IBusCachedPlugin_injectionPort_payload <= debug_bus_cmd_payload_data;
  switch_DebugPlugin_l267 <= pkg_extract(debug_bus_cmd_payload_address,7,2);
  when_DebugPlugin_l271 <= pkg_extract(debug_bus_cmd_payload_data,16);
  when_DebugPlugin_l271_1 <= pkg_extract(debug_bus_cmd_payload_data,24);
  when_DebugPlugin_l272 <= pkg_extract(debug_bus_cmd_payload_data,17);
  when_DebugPlugin_l272_1 <= pkg_extract(debug_bus_cmd_payload_data,25);
  when_DebugPlugin_l273 <= pkg_extract(debug_bus_cmd_payload_data,25);
  when_DebugPlugin_l274 <= pkg_extract(debug_bus_cmd_payload_data,25);
  when_DebugPlugin_l275 <= pkg_extract(debug_bus_cmd_payload_data,18);
  when_DebugPlugin_l275_1 <= pkg_extract(debug_bus_cmd_payload_data,26);
  when_DebugPlugin_l295 <= (execute_arbitration_isValid and execute_DO_EBREAK);
  when_DebugPlugin_l298 <= pkg_toStdLogic(pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_isValid),pkg_toStdLogicVector(memory_arbitration_isValid)) /= pkg_stdLogicVector("00")) = pkg_toStdLogic(false));
  when_DebugPlugin_l311 <= (DebugPlugin_stepIt and IBusCachedPlugin_incomingInstruction);
  debug_resetOut <= DebugPlugin_resetIt_regNext;
  when_DebugPlugin_l327 <= (DebugPlugin_haltIt or DebugPlugin_stepIt);
  when_Pipeline_l124 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_1 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_2 <= ((not writeBack_arbitration_isStuck) and (not CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack));
  when_Pipeline_l124_3 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_4 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_5 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_6 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_7 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_8 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_9 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_10 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_11 <= (not execute_arbitration_isStuck);
  zz_decode_to_execute_SRC1_CTRL_1 <= decode_SRC1_CTRL;
  zz_decode_SRC1_CTRL <= zz_decode_SRC1_CTRL_1;
  when_Pipeline_l124_12 <= (not execute_arbitration_isStuck);
  zz_execute_SRC1_CTRL <= decode_to_execute_SRC1_CTRL;
  when_Pipeline_l124_13 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_14 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_15 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_16 <= (not writeBack_arbitration_isStuck);
  zz_decode_to_execute_ALU_CTRL_1 <= decode_ALU_CTRL;
  zz_decode_ALU_CTRL <= zz_decode_ALU_CTRL_1;
  when_Pipeline_l124_17 <= (not execute_arbitration_isStuck);
  zz_execute_ALU_CTRL <= decode_to_execute_ALU_CTRL;
  zz_decode_to_execute_SRC2_CTRL_1 <= decode_SRC2_CTRL;
  zz_decode_SRC2_CTRL <= zz_decode_SRC2_CTRL_1;
  when_Pipeline_l124_18 <= (not execute_arbitration_isStuck);
  zz_execute_SRC2_CTRL <= decode_to_execute_SRC2_CTRL;
  when_Pipeline_l124_19 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_20 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_21 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_22 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_23 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_24 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_25 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_26 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_27 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_28 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_29 <= (not execute_arbitration_isStuck);
  zz_decode_to_execute_ALU_BITWISE_CTRL_1 <= decode_ALU_BITWISE_CTRL;
  zz_decode_ALU_BITWISE_CTRL <= zz_decode_ALU_BITWISE_CTRL_1;
  when_Pipeline_l124_30 <= (not execute_arbitration_isStuck);
  zz_execute_ALU_BITWISE_CTRL <= decode_to_execute_ALU_BITWISE_CTRL;
  zz_decode_to_execute_SHIFT_CTRL_1 <= decode_SHIFT_CTRL;
  zz_decode_SHIFT_CTRL <= zz_decode_SHIFT_CTRL_1;
  when_Pipeline_l124_31 <= (not execute_arbitration_isStuck);
  zz_execute_SHIFT_CTRL <= decode_to_execute_SHIFT_CTRL;
  when_Pipeline_l124_32 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_33 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_34 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_35 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_36 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_37 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_38 <= (not execute_arbitration_isStuck);
  zz_decode_to_execute_BRANCH_CTRL_1 <= decode_BRANCH_CTRL;
  zz_decode_BRANCH_CTRL <= zz_decode_BRANCH_CTRL_1;
  when_Pipeline_l124_39 <= (not execute_arbitration_isStuck);
  zz_execute_BRANCH_CTRL <= decode_to_execute_BRANCH_CTRL;
  when_Pipeline_l124_40 <= (not execute_arbitration_isStuck);
  zz_decode_to_execute_ENV_CTRL_1 <= decode_ENV_CTRL;
  zz_execute_to_memory_ENV_CTRL_1 <= execute_ENV_CTRL;
  zz_memory_to_writeBack_ENV_CTRL_1 <= memory_ENV_CTRL;
  zz_decode_ENV_CTRL <= zz_decode_ENV_CTRL_1;
  when_Pipeline_l124_41 <= (not execute_arbitration_isStuck);
  zz_execute_ENV_CTRL <= decode_to_execute_ENV_CTRL;
  when_Pipeline_l124_42 <= (not memory_arbitration_isStuck);
  zz_memory_ENV_CTRL <= execute_to_memory_ENV_CTRL;
  when_Pipeline_l124_43 <= (not writeBack_arbitration_isStuck);
  zz_writeBack_ENV_CTRL <= memory_to_writeBack_ENV_CTRL;
  when_Pipeline_l124_44 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_45 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_46 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_47 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_48 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_49 <= (not execute_arbitration_isStuck);
  when_Pipeline_l124_50 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_51 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_52 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_53 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_54 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_55 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_56 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_57 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_58 <= (not writeBack_arbitration_isStuck);
  when_Pipeline_l124_59 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_60 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_61 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_62 <= (not memory_arbitration_isStuck);
  when_Pipeline_l124_63 <= (not writeBack_arbitration_isStuck);
  decode_arbitration_isFlushed <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_flushNext),pkg_cat(pkg_toStdLogicVector(memory_arbitration_flushNext),pkg_toStdLogicVector(execute_arbitration_flushNext))) /= pkg_stdLogicVector("000")) or pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_flushIt),pkg_cat(pkg_toStdLogicVector(memory_arbitration_flushIt),pkg_cat(pkg_toStdLogicVector(execute_arbitration_flushIt),pkg_toStdLogicVector(decode_arbitration_flushIt)))) /= pkg_stdLogicVector("0000")));
  execute_arbitration_isFlushed <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_flushNext),pkg_toStdLogicVector(memory_arbitration_flushNext)) /= pkg_stdLogicVector("00")) or pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_flushIt),pkg_cat(pkg_toStdLogicVector(memory_arbitration_flushIt),pkg_toStdLogicVector(execute_arbitration_flushIt))) /= pkg_stdLogicVector("000")));
  memory_arbitration_isFlushed <= (pkg_toStdLogic(pkg_toStdLogicVector(writeBack_arbitration_flushNext) /= pkg_stdLogicVector("0")) or pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_flushIt),pkg_toStdLogicVector(memory_arbitration_flushIt)) /= pkg_stdLogicVector("00")));
  writeBack_arbitration_isFlushed <= (pkg_toStdLogic(false) or pkg_toStdLogic(pkg_toStdLogicVector(writeBack_arbitration_flushIt) /= pkg_stdLogicVector("0")));
  decode_arbitration_isStuckByOthers <= (decode_arbitration_haltByOther or (((pkg_toStdLogic(false) or execute_arbitration_isStuck) or memory_arbitration_isStuck) or writeBack_arbitration_isStuck));
  decode_arbitration_isStuck <= (decode_arbitration_haltItself or decode_arbitration_isStuckByOthers);
  decode_arbitration_isMoving <= ((not decode_arbitration_isStuck) and (not decode_arbitration_removeIt));
  decode_arbitration_isFiring <= ((decode_arbitration_isValid and (not decode_arbitration_isStuck)) and (not decode_arbitration_removeIt));
  execute_arbitration_isStuckByOthers <= (execute_arbitration_haltByOther or ((pkg_toStdLogic(false) or memory_arbitration_isStuck) or writeBack_arbitration_isStuck));
  execute_arbitration_isStuck <= (execute_arbitration_haltItself or execute_arbitration_isStuckByOthers);
  execute_arbitration_isMoving <= ((not execute_arbitration_isStuck) and (not execute_arbitration_removeIt));
  execute_arbitration_isFiring <= ((execute_arbitration_isValid and (not execute_arbitration_isStuck)) and (not execute_arbitration_removeIt));
  memory_arbitration_isStuckByOthers <= (memory_arbitration_haltByOther or (pkg_toStdLogic(false) or writeBack_arbitration_isStuck));
  memory_arbitration_isStuck <= (memory_arbitration_haltItself or memory_arbitration_isStuckByOthers);
  memory_arbitration_isMoving <= ((not memory_arbitration_isStuck) and (not memory_arbitration_removeIt));
  memory_arbitration_isFiring <= ((memory_arbitration_isValid and (not memory_arbitration_isStuck)) and (not memory_arbitration_removeIt));
  writeBack_arbitration_isStuckByOthers <= (writeBack_arbitration_haltByOther or pkg_toStdLogic(false));
  writeBack_arbitration_isStuck <= (writeBack_arbitration_haltItself or writeBack_arbitration_isStuckByOthers);
  writeBack_arbitration_isMoving <= ((not writeBack_arbitration_isStuck) and (not writeBack_arbitration_removeIt));
  writeBack_arbitration_isFiring <= ((writeBack_arbitration_isValid and (not writeBack_arbitration_isStuck)) and (not writeBack_arbitration_removeIt));
  when_Pipeline_l151 <= ((not execute_arbitration_isStuck) or execute_arbitration_removeIt);
  when_Pipeline_l154 <= ((not decode_arbitration_isStuck) and (not decode_arbitration_removeIt));
  when_Pipeline_l151_1 <= ((not memory_arbitration_isStuck) or memory_arbitration_removeIt);
  when_Pipeline_l154_1 <= ((not execute_arbitration_isStuck) and (not execute_arbitration_removeIt));
  when_Pipeline_l151_2 <= ((not writeBack_arbitration_isStuck) or writeBack_arbitration_removeIt);
  when_Pipeline_l154_2 <= ((not memory_arbitration_isStuck) and (not memory_arbitration_removeIt));
  process(switch_Fetcher_l362)
  begin
    IBusCachedPlugin_injectionPort_ready <= pkg_toStdLogic(false);
    case switch_Fetcher_l362 is
      when "100" =>
        IBusCachedPlugin_injectionPort_ready <= pkg_toStdLogic(true);
      when others =>
    end case;
  end process;

  when_Fetcher_l378 <= (not decode_arbitration_isStuck);
  when_CsrPlugin_l1264 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l1264_1 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l1264_2 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l1264_3 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l1264_4 <= (not execute_arbitration_isStuck);
  when_CsrPlugin_l1264_5 <= (not execute_arbitration_isStuck);
  process(execute_CsrPlugin_csr_768,CsrPlugin_mstatus_MPP,CsrPlugin_mstatus_MPIE,CsrPlugin_mstatus_MIE)
  begin
    zz_CsrPlugin_csrMapping_readDataInit <= pkg_stdLogicVector("00000000000000000000000000000000");
    if execute_CsrPlugin_csr_768 = '1' then
      zz_CsrPlugin_csrMapping_readDataInit(12 downto 11) <= std_logic_vector(CsrPlugin_mstatus_MPP);
      zz_CsrPlugin_csrMapping_readDataInit(7 downto 7) <= pkg_toStdLogicVector(CsrPlugin_mstatus_MPIE);
      zz_CsrPlugin_csrMapping_readDataInit(3 downto 3) <= pkg_toStdLogicVector(CsrPlugin_mstatus_MIE);
    end if;
  end process;

  process(execute_CsrPlugin_csr_836,CsrPlugin_mip_MEIP,CsrPlugin_mip_MTIP,CsrPlugin_mip_MSIP)
  begin
    zz_CsrPlugin_csrMapping_readDataInit_1 <= pkg_stdLogicVector("00000000000000000000000000000000");
    if execute_CsrPlugin_csr_836 = '1' then
      zz_CsrPlugin_csrMapping_readDataInit_1(11 downto 11) <= pkg_toStdLogicVector(CsrPlugin_mip_MEIP);
      zz_CsrPlugin_csrMapping_readDataInit_1(7 downto 7) <= pkg_toStdLogicVector(CsrPlugin_mip_MTIP);
      zz_CsrPlugin_csrMapping_readDataInit_1(3 downto 3) <= pkg_toStdLogicVector(CsrPlugin_mip_MSIP);
    end if;
  end process;

  process(execute_CsrPlugin_csr_772,CsrPlugin_mie_MEIE,CsrPlugin_mie_MTIE,CsrPlugin_mie_MSIE)
  begin
    zz_CsrPlugin_csrMapping_readDataInit_2 <= pkg_stdLogicVector("00000000000000000000000000000000");
    if execute_CsrPlugin_csr_772 = '1' then
      zz_CsrPlugin_csrMapping_readDataInit_2(11 downto 11) <= pkg_toStdLogicVector(CsrPlugin_mie_MEIE);
      zz_CsrPlugin_csrMapping_readDataInit_2(7 downto 7) <= pkg_toStdLogicVector(CsrPlugin_mie_MTIE);
      zz_CsrPlugin_csrMapping_readDataInit_2(3 downto 3) <= pkg_toStdLogicVector(CsrPlugin_mie_MSIE);
    end if;
  end process;

  process(execute_CsrPlugin_csr_833,CsrPlugin_mepc)
  begin
    zz_CsrPlugin_csrMapping_readDataInit_3 <= pkg_stdLogicVector("00000000000000000000000000000000");
    if execute_CsrPlugin_csr_833 = '1' then
      zz_CsrPlugin_csrMapping_readDataInit_3(31 downto 0) <= std_logic_vector(CsrPlugin_mepc);
    end if;
  end process;

  process(execute_CsrPlugin_csr_834,CsrPlugin_mcause_interrupt,CsrPlugin_mcause_exceptionCode)
  begin
    zz_CsrPlugin_csrMapping_readDataInit_4 <= pkg_stdLogicVector("00000000000000000000000000000000");
    if execute_CsrPlugin_csr_834 = '1' then
      zz_CsrPlugin_csrMapping_readDataInit_4(31 downto 31) <= pkg_toStdLogicVector(CsrPlugin_mcause_interrupt);
      zz_CsrPlugin_csrMapping_readDataInit_4(3 downto 0) <= std_logic_vector(CsrPlugin_mcause_exceptionCode);
    end if;
  end process;

  process(execute_CsrPlugin_csr_835,CsrPlugin_mtval)
  begin
    zz_CsrPlugin_csrMapping_readDataInit_5 <= pkg_stdLogicVector("00000000000000000000000000000000");
    if execute_CsrPlugin_csr_835 = '1' then
      zz_CsrPlugin_csrMapping_readDataInit_5(31 downto 0) <= std_logic_vector(CsrPlugin_mtval);
    end if;
  end process;

  CsrPlugin_csrMapping_readDataInit <= (((zz_CsrPlugin_csrMapping_readDataInit or zz_CsrPlugin_csrMapping_readDataInit_1) or (zz_CsrPlugin_csrMapping_readDataInit_2 or zz_CsrPlugin_csrMapping_readDataInit_3)) or (zz_CsrPlugin_csrMapping_readDataInit_4 or zz_CsrPlugin_csrMapping_readDataInit_5));
  when_CsrPlugin_l1297 <= pkg_toStdLogic(CsrPlugin_privilege < unsigned(pkg_extract(execute_CsrPlugin_csrAddress,9,8)));
  when_CsrPlugin_l1302 <= ((not execute_arbitration_isValid) or (not execute_IS_CSR));
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      IBusCachedPlugin_fetchPc_pcReg <= pkg_unsigned("10000000000000000000000000000000");
      IBusCachedPlugin_fetchPc_correctionReg <= pkg_toStdLogic(false);
      IBusCachedPlugin_fetchPc_booted <= pkg_toStdLogic(false);
      IBusCachedPlugin_fetchPc_inc <= pkg_toStdLogic(false);
      zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid <= pkg_toStdLogic(false);
      zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= pkg_toStdLogic(false);
      IBusCachedPlugin_injector_nextPcCalc_valids_0 <= pkg_toStdLogic(false);
      IBusCachedPlugin_injector_nextPcCalc_valids_1 <= pkg_toStdLogic(false);
      IBusCachedPlugin_injector_nextPcCalc_valids_2 <= pkg_toStdLogic(false);
      IBusCachedPlugin_injector_nextPcCalc_valids_3 <= pkg_toStdLogic(false);
      IBusCachedPlugin_injector_nextPcCalc_valids_4 <= pkg_toStdLogic(false);
      IBusCachedPlugin_rspCounter <= zz_IBusCachedPlugin_rspCounter;
      IBusCachedPlugin_rspCounter <= pkg_unsigned("00000000000000000000000000000000");
      DBusCachedPlugin_rspCounter <= zz_DBusCachedPlugin_rspCounter;
      DBusCachedPlugin_rspCounter <= pkg_unsigned("00000000000000000000000000000000");
      zz_3 <= pkg_toStdLogic(true);
      memory_DivPlugin_div_counter_value <= pkg_unsigned("000000");
      HazardSimplePlugin_writeBackBuffer_valid <= pkg_toStdLogic(false);
      CsrPlugin_mstatus_MIE <= pkg_toStdLogic(false);
      CsrPlugin_mstatus_MPIE <= pkg_toStdLogic(false);
      CsrPlugin_mstatus_MPP <= pkg_unsigned("11");
      CsrPlugin_mie_MEIE <= pkg_toStdLogic(false);
      CsrPlugin_mie_MTIE <= pkg_toStdLogic(false);
      CsrPlugin_mie_MSIE <= pkg_toStdLogic(false);
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= pkg_toStdLogic(false);
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= pkg_toStdLogic(false);
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= pkg_toStdLogic(false);
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= pkg_toStdLogic(false);
      CsrPlugin_interrupt_valid <= pkg_toStdLogic(false);
      CsrPlugin_pipelineLiberator_pcValids_0 <= pkg_toStdLogic(false);
      CsrPlugin_pipelineLiberator_pcValids_1 <= pkg_toStdLogic(false);
      CsrPlugin_pipelineLiberator_pcValids_2 <= pkg_toStdLogic(false);
      CsrPlugin_hadException <= pkg_toStdLogic(false);
      execute_CsrPlugin_wfiWake <= pkg_toStdLogic(false);
      execute_arbitration_isValid <= pkg_toStdLogic(false);
      memory_arbitration_isValid <= pkg_toStdLogic(false);
      writeBack_arbitration_isValid <= pkg_toStdLogic(false);
      switch_Fetcher_l362 <= pkg_unsigned("000");
    elsif rising_edge(io_mainClk) then
      if IBusCachedPlugin_fetchPc_correction = '1' then
        IBusCachedPlugin_fetchPc_correctionReg <= pkg_toStdLogic(true);
      end if;
      if IBusCachedPlugin_fetchPc_output_fire = '1' then
        IBusCachedPlugin_fetchPc_correctionReg <= pkg_toStdLogic(false);
      end if;
      IBusCachedPlugin_fetchPc_booted <= pkg_toStdLogic(true);
      if when_Fetcher_l131 = '1' then
        IBusCachedPlugin_fetchPc_inc <= pkg_toStdLogic(false);
      end if;
      if IBusCachedPlugin_fetchPc_output_fire_1 = '1' then
        IBusCachedPlugin_fetchPc_inc <= pkg_toStdLogic(true);
      end if;
      if when_Fetcher_l131_1 = '1' then
        IBusCachedPlugin_fetchPc_inc <= pkg_toStdLogic(false);
      end if;
      if when_Fetcher_l158 = '1' then
        IBusCachedPlugin_fetchPc_pcReg <= IBusCachedPlugin_fetchPc_pc;
      end if;
      if IBusCachedPlugin_iBusRsp_flush = '1' then
        zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid <= pkg_toStdLogic(false);
      end if;
      if IBusCachedPlugin_iBusRsp_stages_0_output_ready = '1' then
        zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_0_output_valid and (not pkg_toStdLogic(false)));
      end if;
      if IBusCachedPlugin_iBusRsp_flush = '1' then
        zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= pkg_toStdLogic(false);
      end if;
      if IBusCachedPlugin_iBusRsp_stages_1_output_ready = '1' then
        zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_1_output_valid and (not IBusCachedPlugin_iBusRsp_flush));
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= pkg_toStdLogic(false);
      end if;
      if when_Fetcher_l329 = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= pkg_toStdLogic(true);
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= pkg_toStdLogic(false);
      end if;
      if when_Fetcher_l329_1 = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_0;
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= pkg_toStdLogic(false);
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= pkg_toStdLogic(false);
      end if;
      if when_Fetcher_l329_2 = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= pkg_toStdLogic(false);
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= pkg_toStdLogic(false);
      end if;
      if when_Fetcher_l329_3 = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= pkg_toStdLogic(false);
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= pkg_toStdLogic(false);
      end if;
      if when_Fetcher_l329_4 = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= IBusCachedPlugin_injector_nextPcCalc_valids_3;
      end if;
      if IBusCachedPlugin_fetchPc_flushed = '1' then
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= pkg_toStdLogic(false);
      end if;
      if iBus_rsp_valid = '1' then
        IBusCachedPlugin_rspCounter <= (IBusCachedPlugin_rspCounter + pkg_unsigned("00000000000000000000000000000001"));
      end if;
      if dBus_rsp_valid = '1' then
        DBusCachedPlugin_rspCounter <= (DBusCachedPlugin_rspCounter + pkg_unsigned("00000000000000000000000000000001"));
      end if;
      zz_3 <= pkg_toStdLogic(false);
      memory_DivPlugin_div_counter_value <= memory_DivPlugin_div_counter_valueNext;
      HazardSimplePlugin_writeBackBuffer_valid <= HazardSimplePlugin_writeBackWrites_valid;
      if when_CsrPlugin_l909 = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= pkg_toStdLogic(false);
      else
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
      end if;
      if when_CsrPlugin_l909_1 = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= (CsrPlugin_exceptionPortCtrl_exceptionValids_decode and (not decode_arbitration_isStuck));
      else
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
      end if;
      if when_CsrPlugin_l909_2 = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= (CsrPlugin_exceptionPortCtrl_exceptionValids_execute and (not execute_arbitration_isStuck));
      else
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
      end if;
      if when_CsrPlugin_l909_3 = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= (CsrPlugin_exceptionPortCtrl_exceptionValids_memory and (not memory_arbitration_isStuck));
      else
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= pkg_toStdLogic(false);
      end if;
      CsrPlugin_interrupt_valid <= pkg_toStdLogic(false);
      if when_CsrPlugin_l946 = '1' then
        if when_CsrPlugin_l952 = '1' then
          CsrPlugin_interrupt_valid <= pkg_toStdLogic(true);
        end if;
        if when_CsrPlugin_l952_1 = '1' then
          CsrPlugin_interrupt_valid <= pkg_toStdLogic(true);
        end if;
        if when_CsrPlugin_l952_2 = '1' then
          CsrPlugin_interrupt_valid <= pkg_toStdLogic(true);
        end if;
      end if;
      if CsrPlugin_pipelineLiberator_active = '1' then
        if when_CsrPlugin_l980 = '1' then
          CsrPlugin_pipelineLiberator_pcValids_0 <= pkg_toStdLogic(true);
        end if;
        if when_CsrPlugin_l980_1 = '1' then
          CsrPlugin_pipelineLiberator_pcValids_1 <= CsrPlugin_pipelineLiberator_pcValids_0;
        end if;
        if when_CsrPlugin_l980_2 = '1' then
          CsrPlugin_pipelineLiberator_pcValids_2 <= CsrPlugin_pipelineLiberator_pcValids_1;
        end if;
      end if;
      if when_CsrPlugin_l985 = '1' then
        CsrPlugin_pipelineLiberator_pcValids_0 <= pkg_toStdLogic(false);
        CsrPlugin_pipelineLiberator_pcValids_1 <= pkg_toStdLogic(false);
        CsrPlugin_pipelineLiberator_pcValids_2 <= pkg_toStdLogic(false);
      end if;
      if CsrPlugin_interruptJump = '1' then
        CsrPlugin_interrupt_valid <= pkg_toStdLogic(false);
      end if;
      CsrPlugin_hadException <= CsrPlugin_exception;
      if when_CsrPlugin_l1019 = '1' then
        case CsrPlugin_targetPrivilege is
          when "11" =>
            CsrPlugin_mstatus_MIE <= pkg_toStdLogic(false);
            CsrPlugin_mstatus_MPIE <= CsrPlugin_mstatus_MIE;
            CsrPlugin_mstatus_MPP <= CsrPlugin_privilege;
          when others =>
        end case;
      end if;
      if when_CsrPlugin_l1064 = '1' then
        case switch_CsrPlugin_l1068 is
          when "11" =>
            CsrPlugin_mstatus_MPP <= pkg_unsigned("00");
            CsrPlugin_mstatus_MIE <= CsrPlugin_mstatus_MPIE;
            CsrPlugin_mstatus_MPIE <= pkg_toStdLogic(true);
          when others =>
        end case;
      end if;
      execute_CsrPlugin_wfiWake <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(zz_when_CsrPlugin_l952_2),pkg_cat(pkg_toStdLogicVector(zz_when_CsrPlugin_l952_1),pkg_toStdLogicVector(zz_when_CsrPlugin_l952))) /= pkg_stdLogicVector("000")) or CsrPlugin_thirdPartyWake);
      if when_Pipeline_l151 = '1' then
        execute_arbitration_isValid <= pkg_toStdLogic(false);
      end if;
      if when_Pipeline_l154 = '1' then
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end if;
      if when_Pipeline_l151_1 = '1' then
        memory_arbitration_isValid <= pkg_toStdLogic(false);
      end if;
      if when_Pipeline_l154_1 = '1' then
        memory_arbitration_isValid <= execute_arbitration_isValid;
      end if;
      if when_Pipeline_l151_2 = '1' then
        writeBack_arbitration_isValid <= pkg_toStdLogic(false);
      end if;
      if when_Pipeline_l154_2 = '1' then
        writeBack_arbitration_isValid <= memory_arbitration_isValid;
      end if;
      case switch_Fetcher_l362 is
        when "000" =>
          if IBusCachedPlugin_injectionPort_valid = '1' then
            switch_Fetcher_l362 <= pkg_unsigned("001");
          end if;
        when "001" =>
          switch_Fetcher_l362 <= pkg_unsigned("010");
        when "010" =>
          switch_Fetcher_l362 <= pkg_unsigned("011");
        when "011" =>
          if when_Fetcher_l378 = '1' then
            switch_Fetcher_l362 <= pkg_unsigned("100");
          end if;
        when "100" =>
          switch_Fetcher_l362 <= pkg_unsigned("000");
        when others =>
      end case;
      if execute_CsrPlugin_csr_768 = '1' then
        if execute_CsrPlugin_writeEnable = '1' then
          CsrPlugin_mstatus_MPP <= unsigned(pkg_extract(CsrPlugin_csrMapping_writeDataSignal,12,11));
          CsrPlugin_mstatus_MPIE <= pkg_extract(CsrPlugin_csrMapping_writeDataSignal,7);
          CsrPlugin_mstatus_MIE <= pkg_extract(CsrPlugin_csrMapping_writeDataSignal,3);
        end if;
      end if;
      if execute_CsrPlugin_csr_772 = '1' then
        if execute_CsrPlugin_writeEnable = '1' then
          CsrPlugin_mie_MEIE <= pkg_extract(CsrPlugin_csrMapping_writeDataSignal,11);
          CsrPlugin_mie_MTIE <= pkg_extract(CsrPlugin_csrMapping_writeDataSignal,7);
          CsrPlugin_mie_MSIE <= pkg_extract(CsrPlugin_csrMapping_writeDataSignal,3);
        end if;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if IBusCachedPlugin_iBusRsp_stages_0_output_ready = '1' then
        zz_IBusCachedPlugin_iBusRsp_stages_0_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_0_output_payload;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_1_output_ready = '1' then
        zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_payload;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_0_output_ready = '1' then
        IBusCachedPlugin_predictor_writeLast_valid <= IBusCachedPlugin_predictor_historyWriteDelayPatched_valid;
        IBusCachedPlugin_predictor_writeLast_payload_address <= IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_address;
        IBusCachedPlugin_predictor_writeLast_payload_data_source <= IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_source;
        IBusCachedPlugin_predictor_writeLast_payload_data_branchWish <= IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_branchWish;
        IBusCachedPlugin_predictor_writeLast_payload_data_target <= IBusCachedPlugin_predictor_historyWriteDelayPatched_payload_data_target;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_0_input_ready = '1' then
        IBusCachedPlugin_predictor_buffer_pcCorrected <= IBusCachedPlugin_fetchPc_corrected;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_0_output_ready = '1' then
        IBusCachedPlugin_predictor_line_source <= IBusCachedPlugin_predictor_buffer_line_source;
        IBusCachedPlugin_predictor_line_branchWish <= IBusCachedPlugin_predictor_buffer_line_branchWish;
        IBusCachedPlugin_predictor_line_target <= IBusCachedPlugin_predictor_buffer_line_target;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_0_output_ready = '1' then
        IBusCachedPlugin_predictor_buffer_hazard_regNextWhen <= IBusCachedPlugin_predictor_buffer_hazard;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_1_output_ready = '1' then
        IBusCachedPlugin_predictor_iBusRspContext_hazard <= IBusCachedPlugin_predictor_fetchContext_hazard;
        IBusCachedPlugin_predictor_iBusRspContext_hit <= IBusCachedPlugin_predictor_fetchContext_hit;
        IBusCachedPlugin_predictor_iBusRspContext_line_source <= IBusCachedPlugin_predictor_fetchContext_line_source;
        IBusCachedPlugin_predictor_iBusRspContext_line_branchWish <= IBusCachedPlugin_predictor_fetchContext_line_branchWish;
        IBusCachedPlugin_predictor_iBusRspContext_line_target <= IBusCachedPlugin_predictor_fetchContext_line_target;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_1_input_ready = '1' then
        IBusCachedPlugin_s1_tightlyCoupledHit <= IBusCachedPlugin_s0_tightlyCoupledHit;
      end if;
      if IBusCachedPlugin_iBusRsp_stages_2_input_ready = '1' then
        IBusCachedPlugin_s2_tightlyCoupledHit <= IBusCachedPlugin_s1_tightlyCoupledHit;
      end if;
      if when_MulDivIterativePlugin_l126 = '1' then
        memory_DivPlugin_div_done <= pkg_toStdLogic(true);
      end if;
      if when_MulDivIterativePlugin_l126_1 = '1' then
        memory_DivPlugin_div_done <= pkg_toStdLogic(false);
      end if;
      if when_MulDivIterativePlugin_l128 = '1' then
        if when_MulDivIterativePlugin_l132 = '1' then
          memory_DivPlugin_rs1(31 downto 0) <= memory_DivPlugin_div_stage_0_outNumerator;
          memory_DivPlugin_accumulator(31 downto 0) <= memory_DivPlugin_div_stage_0_outRemainder;
          if when_MulDivIterativePlugin_l151 = '1' then
            memory_DivPlugin_div_result <= pkg_resize(std_logic_vector(signed((unsigned(pkg_cat(pkg_toStdLogicVector(memory_DivPlugin_div_needRevert),std_logic_vector(pkg_mux(memory_DivPlugin_div_needRevert,pkg_not(zz_memory_DivPlugin_div_result),zz_memory_DivPlugin_div_result)))) + pkg_resize(unsigned(pkg_toStdLogicVector(memory_DivPlugin_div_needRevert)),33)))),32);
          end if;
        end if;
      end if;
      if when_MulDivIterativePlugin_l162 = '1' then
        memory_DivPlugin_accumulator <= pkg_unsigned("00000000000000000000000000000000000000000000000000000000000000000");
        memory_DivPlugin_rs1 <= (unsigned(pkg_mux(zz_memory_DivPlugin_rs1,pkg_not(zz_memory_DivPlugin_rs1_1),zz_memory_DivPlugin_rs1_1)) + pkg_resize(unsigned(pkg_toStdLogicVector(zz_memory_DivPlugin_rs1)),33));
        memory_DivPlugin_rs2 <= (unsigned(pkg_mux(zz_memory_DivPlugin_rs2,pkg_not(execute_RS2),execute_RS2)) + pkg_resize(unsigned(pkg_toStdLogicVector(zz_memory_DivPlugin_rs2)),32));
        memory_DivPlugin_div_needRevert <= ((zz_memory_DivPlugin_rs1 xor (zz_memory_DivPlugin_rs2 and (not pkg_extract(execute_INSTRUCTION,13)))) and (not ((pkg_toStdLogic(execute_RS2 = pkg_stdLogicVector("00000000000000000000000000000000")) and execute_IS_RS2_SIGNED) and (not pkg_extract(execute_INSTRUCTION,13)))));
      end if;
      HazardSimplePlugin_writeBackBuffer_payload_address <= HazardSimplePlugin_writeBackWrites_payload_address;
      HazardSimplePlugin_writeBackBuffer_payload_data <= HazardSimplePlugin_writeBackWrites_payload_data;
      CsrPlugin_mip_MEIP <= externalInterrupt;
      CsrPlugin_mip_MTIP <= timerInterrupt;
      CsrPlugin_mip_MSIP <= softwareInterrupt;
      CsrPlugin_mcycle <= (CsrPlugin_mcycle + pkg_unsigned("0000000000000000000000000000000000000000000000000000000000000001"));
      if writeBack_arbitration_isFiring = '1' then
        CsrPlugin_minstret <= (CsrPlugin_minstret + pkg_unsigned("0000000000000000000000000000000000000000000000000000000000000001"));
      end if;
      if zz_when = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionContext_code <= pkg_mux(zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1,IBusCachedPlugin_decodeExceptionPort_payload_code,decodeExceptionPort_payload_code);
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= pkg_mux(zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1,IBusCachedPlugin_decodeExceptionPort_payload_badAddr,decodeExceptionPort_payload_badAddr);
      end if;
      if BranchPlugin_branchExceptionPort_valid = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionContext_code <= BranchPlugin_branchExceptionPort_payload_code;
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= BranchPlugin_branchExceptionPort_payload_badAddr;
      end if;
      if DBusCachedPlugin_exceptionBus_valid = '1' then
        CsrPlugin_exceptionPortCtrl_exceptionContext_code <= DBusCachedPlugin_exceptionBus_payload_code;
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= DBusCachedPlugin_exceptionBus_payload_badAddr;
      end if;
      if when_CsrPlugin_l946 = '1' then
        if when_CsrPlugin_l952 = '1' then
          CsrPlugin_interrupt_code <= pkg_unsigned("0111");
          CsrPlugin_interrupt_targetPrivilege <= pkg_unsigned("11");
        end if;
        if when_CsrPlugin_l952_1 = '1' then
          CsrPlugin_interrupt_code <= pkg_unsigned("0011");
          CsrPlugin_interrupt_targetPrivilege <= pkg_unsigned("11");
        end if;
        if when_CsrPlugin_l952_2 = '1' then
          CsrPlugin_interrupt_code <= pkg_unsigned("1011");
          CsrPlugin_interrupt_targetPrivilege <= pkg_unsigned("11");
        end if;
      end if;
      if when_CsrPlugin_l1019 = '1' then
        case CsrPlugin_targetPrivilege is
          when "11" =>
            CsrPlugin_mcause_interrupt <= (not CsrPlugin_hadException);
            CsrPlugin_mcause_exceptionCode <= CsrPlugin_trapCause;
            CsrPlugin_mepc <= writeBack_PC;
            if CsrPlugin_hadException = '1' then
              CsrPlugin_mtval <= CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
            end if;
          when others =>
        end case;
      end if;
      if when_Pipeline_l124 = '1' then
        decode_to_execute_PC <= decode_PC;
      end if;
      if when_Pipeline_l124_1 = '1' then
        execute_to_memory_PC <= zz_execute_SRC2;
      end if;
      if when_Pipeline_l124_2 = '1' then
        memory_to_writeBack_PC <= memory_PC;
      end if;
      if when_Pipeline_l124_3 = '1' then
        decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
      end if;
      if when_Pipeline_l124_4 = '1' then
        execute_to_memory_INSTRUCTION <= execute_INSTRUCTION;
      end if;
      if when_Pipeline_l124_5 = '1' then
        memory_to_writeBack_INSTRUCTION <= memory_INSTRUCTION;
      end if;
      if when_Pipeline_l124_6 = '1' then
        decode_to_execute_FORMAL_PC_NEXT <= decode_FORMAL_PC_NEXT;
      end if;
      if when_Pipeline_l124_7 = '1' then
        execute_to_memory_FORMAL_PC_NEXT <= execute_FORMAL_PC_NEXT;
      end if;
      if when_Pipeline_l124_8 = '1' then
        memory_to_writeBack_FORMAL_PC_NEXT <= zz_memory_to_writeBack_FORMAL_PC_NEXT;
      end if;
      if when_Pipeline_l124_9 = '1' then
        decode_to_execute_PREDICTION_CONTEXT_hazard <= decode_PREDICTION_CONTEXT_hazard;
        decode_to_execute_PREDICTION_CONTEXT_hit <= decode_PREDICTION_CONTEXT_hit;
        decode_to_execute_PREDICTION_CONTEXT_line_source <= decode_PREDICTION_CONTEXT_line_source;
        decode_to_execute_PREDICTION_CONTEXT_line_branchWish <= decode_PREDICTION_CONTEXT_line_branchWish;
        decode_to_execute_PREDICTION_CONTEXT_line_target <= decode_PREDICTION_CONTEXT_line_target;
      end if;
      if when_Pipeline_l124_10 = '1' then
        execute_to_memory_PREDICTION_CONTEXT_hazard <= execute_PREDICTION_CONTEXT_hazard;
        execute_to_memory_PREDICTION_CONTEXT_hit <= execute_PREDICTION_CONTEXT_hit;
        execute_to_memory_PREDICTION_CONTEXT_line_source <= execute_PREDICTION_CONTEXT_line_source;
        execute_to_memory_PREDICTION_CONTEXT_line_branchWish <= execute_PREDICTION_CONTEXT_line_branchWish;
        execute_to_memory_PREDICTION_CONTEXT_line_target <= execute_PREDICTION_CONTEXT_line_target;
      end if;
      if when_Pipeline_l124_11 = '1' then
        decode_to_execute_MEMORY_FORCE_CONSTISTENCY <= decode_MEMORY_FORCE_CONSTISTENCY;
      end if;
      if when_Pipeline_l124_12 = '1' then
        decode_to_execute_SRC1_CTRL <= zz_decode_to_execute_SRC1_CTRL;
      end if;
      if when_Pipeline_l124_13 = '1' then
        decode_to_execute_SRC_USE_SUB_LESS <= decode_SRC_USE_SUB_LESS;
      end if;
      if when_Pipeline_l124_14 = '1' then
        decode_to_execute_MEMORY_ENABLE <= decode_MEMORY_ENABLE;
      end if;
      if when_Pipeline_l124_15 = '1' then
        execute_to_memory_MEMORY_ENABLE <= execute_MEMORY_ENABLE;
      end if;
      if when_Pipeline_l124_16 = '1' then
        memory_to_writeBack_MEMORY_ENABLE <= memory_MEMORY_ENABLE;
      end if;
      if when_Pipeline_l124_17 = '1' then
        decode_to_execute_ALU_CTRL <= zz_decode_to_execute_ALU_CTRL;
      end if;
      if when_Pipeline_l124_18 = '1' then
        decode_to_execute_SRC2_CTRL <= zz_decode_to_execute_SRC2_CTRL;
      end if;
      if when_Pipeline_l124_19 = '1' then
        decode_to_execute_REGFILE_WRITE_VALID <= decode_REGFILE_WRITE_VALID;
      end if;
      if when_Pipeline_l124_20 = '1' then
        execute_to_memory_REGFILE_WRITE_VALID <= execute_REGFILE_WRITE_VALID;
      end if;
      if when_Pipeline_l124_21 = '1' then
        memory_to_writeBack_REGFILE_WRITE_VALID <= memory_REGFILE_WRITE_VALID;
      end if;
      if when_Pipeline_l124_22 = '1' then
        decode_to_execute_BYPASSABLE_EXECUTE_STAGE <= decode_BYPASSABLE_EXECUTE_STAGE;
      end if;
      if when_Pipeline_l124_23 = '1' then
        decode_to_execute_BYPASSABLE_MEMORY_STAGE <= decode_BYPASSABLE_MEMORY_STAGE;
      end if;
      if when_Pipeline_l124_24 = '1' then
        execute_to_memory_BYPASSABLE_MEMORY_STAGE <= execute_BYPASSABLE_MEMORY_STAGE;
      end if;
      if when_Pipeline_l124_25 = '1' then
        decode_to_execute_MEMORY_WR <= decode_MEMORY_WR;
      end if;
      if when_Pipeline_l124_26 = '1' then
        execute_to_memory_MEMORY_WR <= execute_MEMORY_WR;
      end if;
      if when_Pipeline_l124_27 = '1' then
        memory_to_writeBack_MEMORY_WR <= memory_MEMORY_WR;
      end if;
      if when_Pipeline_l124_28 = '1' then
        decode_to_execute_MEMORY_MANAGMENT <= decode_MEMORY_MANAGMENT;
      end if;
      if when_Pipeline_l124_29 = '1' then
        decode_to_execute_SRC_LESS_UNSIGNED <= decode_SRC_LESS_UNSIGNED;
      end if;
      if when_Pipeline_l124_30 = '1' then
        decode_to_execute_ALU_BITWISE_CTRL <= zz_decode_to_execute_ALU_BITWISE_CTRL;
      end if;
      if when_Pipeline_l124_31 = '1' then
        decode_to_execute_SHIFT_CTRL <= zz_decode_to_execute_SHIFT_CTRL;
      end if;
      if when_Pipeline_l124_32 = '1' then
        decode_to_execute_IS_MUL <= decode_IS_MUL;
      end if;
      if when_Pipeline_l124_33 = '1' then
        execute_to_memory_IS_MUL <= execute_IS_MUL;
      end if;
      if when_Pipeline_l124_34 = '1' then
        memory_to_writeBack_IS_MUL <= memory_IS_MUL;
      end if;
      if when_Pipeline_l124_35 = '1' then
        decode_to_execute_IS_DIV <= decode_IS_DIV;
      end if;
      if when_Pipeline_l124_36 = '1' then
        execute_to_memory_IS_DIV <= execute_IS_DIV;
      end if;
      if when_Pipeline_l124_37 = '1' then
        decode_to_execute_IS_RS1_SIGNED <= decode_IS_RS1_SIGNED;
      end if;
      if when_Pipeline_l124_38 = '1' then
        decode_to_execute_IS_RS2_SIGNED <= decode_IS_RS2_SIGNED;
      end if;
      if when_Pipeline_l124_39 = '1' then
        decode_to_execute_BRANCH_CTRL <= zz_decode_to_execute_BRANCH_CTRL;
      end if;
      if when_Pipeline_l124_40 = '1' then
        decode_to_execute_IS_CSR <= decode_IS_CSR;
      end if;
      if when_Pipeline_l124_41 = '1' then
        decode_to_execute_ENV_CTRL <= zz_decode_to_execute_ENV_CTRL;
      end if;
      if when_Pipeline_l124_42 = '1' then
        execute_to_memory_ENV_CTRL <= zz_execute_to_memory_ENV_CTRL;
      end if;
      if when_Pipeline_l124_43 = '1' then
        memory_to_writeBack_ENV_CTRL <= zz_memory_to_writeBack_ENV_CTRL;
      end if;
      if when_Pipeline_l124_44 = '1' then
        decode_to_execute_RS1 <= decode_RS1;
      end if;
      if when_Pipeline_l124_45 = '1' then
        decode_to_execute_RS2 <= decode_RS2;
      end if;
      if when_Pipeline_l124_46 = '1' then
        decode_to_execute_SRC2_FORCE_ZERO <= decode_SRC2_FORCE_ZERO;
      end if;
      if when_Pipeline_l124_47 = '1' then
        decode_to_execute_CSR_WRITE_OPCODE <= decode_CSR_WRITE_OPCODE;
      end if;
      if when_Pipeline_l124_48 = '1' then
        decode_to_execute_CSR_READ_OPCODE <= decode_CSR_READ_OPCODE;
      end if;
      if when_Pipeline_l124_49 = '1' then
        decode_to_execute_DO_EBREAK <= decode_DO_EBREAK;
      end if;
      if when_Pipeline_l124_50 = '1' then
        execute_to_memory_MEMORY_STORE_DATA_RF <= execute_MEMORY_STORE_DATA_RF;
      end if;
      if when_Pipeline_l124_51 = '1' then
        memory_to_writeBack_MEMORY_STORE_DATA_RF <= memory_MEMORY_STORE_DATA_RF;
      end if;
      if when_Pipeline_l124_52 = '1' then
        execute_to_memory_REGFILE_WRITE_DATA <= zz_decode_RS2_1;
      end if;
      if when_Pipeline_l124_53 = '1' then
        memory_to_writeBack_REGFILE_WRITE_DATA <= zz_decode_RS2;
      end if;
      if when_Pipeline_l124_54 = '1' then
        execute_to_memory_MUL_LL <= execute_MUL_LL;
      end if;
      if when_Pipeline_l124_55 = '1' then
        execute_to_memory_MUL_LH <= execute_MUL_LH;
      end if;
      if when_Pipeline_l124_56 = '1' then
        execute_to_memory_MUL_HL <= execute_MUL_HL;
      end if;
      if when_Pipeline_l124_57 = '1' then
        execute_to_memory_MUL_HH <= execute_MUL_HH;
      end if;
      if when_Pipeline_l124_58 = '1' then
        memory_to_writeBack_MUL_HH <= memory_MUL_HH;
      end if;
      if when_Pipeline_l124_59 = '1' then
        execute_to_memory_BRANCH_DO <= execute_BRANCH_DO;
      end if;
      if when_Pipeline_l124_60 = '1' then
        execute_to_memory_BRANCH_CALC <= execute_BRANCH_CALC;
      end if;
      if when_Pipeline_l124_61 = '1' then
        execute_to_memory_NEXT_PC2 <= execute_NEXT_PC2;
      end if;
      if when_Pipeline_l124_62 = '1' then
        execute_to_memory_TARGET_MISSMATCH2 <= execute_TARGET_MISSMATCH2;
      end if;
      if when_Pipeline_l124_63 = '1' then
        memory_to_writeBack_MUL_LOW <= memory_MUL_LOW;
      end if;
      if when_CsrPlugin_l1264 = '1' then
        execute_CsrPlugin_csr_768 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,31,20) = pkg_stdLogicVector("001100000000"));
      end if;
      if when_CsrPlugin_l1264_1 = '1' then
        execute_CsrPlugin_csr_836 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,31,20) = pkg_stdLogicVector("001101000100"));
      end if;
      if when_CsrPlugin_l1264_2 = '1' then
        execute_CsrPlugin_csr_772 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,31,20) = pkg_stdLogicVector("001100000100"));
      end if;
      if when_CsrPlugin_l1264_3 = '1' then
        execute_CsrPlugin_csr_833 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,31,20) = pkg_stdLogicVector("001101000001"));
      end if;
      if when_CsrPlugin_l1264_4 = '1' then
        execute_CsrPlugin_csr_834 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,31,20) = pkg_stdLogicVector("001101000010"));
      end if;
      if when_CsrPlugin_l1264_5 = '1' then
        execute_CsrPlugin_csr_835 <= pkg_toStdLogic(pkg_extract(decode_INSTRUCTION,31,20) = pkg_stdLogicVector("001101000011"));
      end if;
      if execute_CsrPlugin_csr_836 = '1' then
        if execute_CsrPlugin_writeEnable = '1' then
          CsrPlugin_mip_MSIP <= pkg_extract(CsrPlugin_csrMapping_writeDataSignal,3);
        end if;
      end if;
      if execute_CsrPlugin_csr_833 = '1' then
        if execute_CsrPlugin_writeEnable = '1' then
          CsrPlugin_mepc <= unsigned(pkg_extract(CsrPlugin_csrMapping_writeDataSignal,31,0));
        end if;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      DebugPlugin_firstCycle <= pkg_toStdLogic(false);
      if debug_bus_cmd_ready_read_buffer = '1' then
        DebugPlugin_firstCycle <= pkg_toStdLogic(true);
      end if;
      DebugPlugin_secondCycle <= DebugPlugin_firstCycle;
      DebugPlugin_isPipBusy <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(writeBack_arbitration_isValid),pkg_cat(pkg_toStdLogicVector(memory_arbitration_isValid),pkg_cat(pkg_toStdLogicVector(execute_arbitration_isValid),pkg_toStdLogicVector(decode_arbitration_isValid)))) /= pkg_stdLogicVector("0000")) or IBusCachedPlugin_incomingInstruction);
      if writeBack_arbitration_isValid = '1' then
        DebugPlugin_busReadDataReg <= zz_decode_RS2_2;
      end if;
      zz_when_DebugPlugin_l244 <= pkg_extract(debug_bus_cmd_payload_address,2);
      if when_DebugPlugin_l295 = '1' then
        DebugPlugin_busReadDataReg <= std_logic_vector(execute_PC);
      end if;
      DebugPlugin_resetIt_regNext <= DebugPlugin_resetIt;
    end if;
  end process;

  process(io_mainClk, resetCtrl_systemReset)
  begin
    if resetCtrl_systemReset = '1' then
      DebugPlugin_resetIt <= pkg_toStdLogic(false);
      DebugPlugin_haltIt <= pkg_toStdLogic(false);
      DebugPlugin_stepIt <= pkg_toStdLogic(false);
      DebugPlugin_godmode <= pkg_toStdLogic(false);
      DebugPlugin_haltedByBreak <= pkg_toStdLogic(false);
      DebugPlugin_debugUsed <= pkg_toStdLogic(false);
      DebugPlugin_disableEbreak <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if when_DebugPlugin_l225 = '1' then
        DebugPlugin_godmode <= pkg_toStdLogic(true);
      end if;
      if debug_bus_cmd_valid = '1' then
        DebugPlugin_debugUsed <= pkg_toStdLogic(true);
      end if;
      if debug_bus_cmd_valid = '1' then
        case switch_DebugPlugin_l267 is
          when "000000" =>
            if debug_bus_cmd_payload_wr = '1' then
              DebugPlugin_stepIt <= pkg_extract(debug_bus_cmd_payload_data,4);
              if when_DebugPlugin_l271 = '1' then
                DebugPlugin_resetIt <= pkg_toStdLogic(true);
              end if;
              if when_DebugPlugin_l271_1 = '1' then
                DebugPlugin_resetIt <= pkg_toStdLogic(false);
              end if;
              if when_DebugPlugin_l272 = '1' then
                DebugPlugin_haltIt <= pkg_toStdLogic(true);
              end if;
              if when_DebugPlugin_l272_1 = '1' then
                DebugPlugin_haltIt <= pkg_toStdLogic(false);
              end if;
              if when_DebugPlugin_l273 = '1' then
                DebugPlugin_haltedByBreak <= pkg_toStdLogic(false);
              end if;
              if when_DebugPlugin_l274 = '1' then
                DebugPlugin_godmode <= pkg_toStdLogic(false);
              end if;
              if when_DebugPlugin_l275 = '1' then
                DebugPlugin_disableEbreak <= pkg_toStdLogic(true);
              end if;
              if when_DebugPlugin_l275_1 = '1' then
                DebugPlugin_disableEbreak <= pkg_toStdLogic(false);
              end if;
            end if;
          when others =>
        end case;
      end if;
      if when_DebugPlugin_l295 = '1' then
        if when_DebugPlugin_l298 = '1' then
          DebugPlugin_haltIt <= pkg_toStdLogic(true);
          DebugPlugin_haltedByBreak <= pkg_toStdLogic(true);
        end if;
      end if;
      if when_DebugPlugin_l311 = '1' then
        if decode_arbitration_isValid = '1' then
          DebugPlugin_haltIt <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity StreamFork_2 is
  port(
    io_input_valid : in std_logic;
    io_input_ready : out std_logic;
    io_input_payload_wr : in std_logic;
    io_input_payload_uncached : in std_logic;
    io_input_payload_address : in unsigned(31 downto 0);
    io_input_payload_data : in std_logic_vector(31 downto 0);
    io_input_payload_mask : in std_logic_vector(3 downto 0);
    io_input_payload_size : in unsigned(2 downto 0);
    io_input_payload_last : in std_logic;
    io_outputs_0_valid : out std_logic;
    io_outputs_0_ready : in std_logic;
    io_outputs_0_payload_wr : out std_logic;
    io_outputs_0_payload_uncached : out std_logic;
    io_outputs_0_payload_address : out unsigned(31 downto 0);
    io_outputs_0_payload_data : out std_logic_vector(31 downto 0);
    io_outputs_0_payload_mask : out std_logic_vector(3 downto 0);
    io_outputs_0_payload_size : out unsigned(2 downto 0);
    io_outputs_0_payload_last : out std_logic;
    io_outputs_1_valid : out std_logic;
    io_outputs_1_ready : in std_logic;
    io_outputs_1_payload_wr : out std_logic;
    io_outputs_1_payload_uncached : out std_logic;
    io_outputs_1_payload_address : out unsigned(31 downto 0);
    io_outputs_1_payload_data : out std_logic_vector(31 downto 0);
    io_outputs_1_payload_mask : out std_logic_vector(3 downto 0);
    io_outputs_1_payload_size : out unsigned(2 downto 0);
    io_outputs_1_payload_last : out std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end StreamFork_2;

architecture arch of StreamFork_2 is
  signal io_outputs_0_valid_read_buffer : std_logic;
  signal io_outputs_1_valid_read_buffer : std_logic;
  signal io_input_ready_read_buffer : std_logic;

  signal zz_io_outputs_0_valid : std_logic;
  signal zz_io_outputs_1_valid : std_logic;
  signal when_Stream_l817 : std_logic;
  signal when_Stream_l817_1 : std_logic;
  signal io_outputs_0_fire : std_logic;
  signal io_outputs_1_fire : std_logic;
begin
  io_outputs_0_valid <= io_outputs_0_valid_read_buffer;
  io_outputs_1_valid <= io_outputs_1_valid_read_buffer;
  io_input_ready <= io_input_ready_read_buffer;
  process(when_Stream_l817,when_Stream_l817_1)
  begin
    io_input_ready_read_buffer <= pkg_toStdLogic(true);
    if when_Stream_l817 = '1' then
      io_input_ready_read_buffer <= pkg_toStdLogic(false);
    end if;
    if when_Stream_l817_1 = '1' then
      io_input_ready_read_buffer <= pkg_toStdLogic(false);
    end if;
  end process;

  when_Stream_l817 <= ((not io_outputs_0_ready) and zz_io_outputs_0_valid);
  when_Stream_l817_1 <= ((not io_outputs_1_ready) and zz_io_outputs_1_valid);
  io_outputs_0_valid_read_buffer <= (io_input_valid and zz_io_outputs_0_valid);
  io_outputs_0_payload_wr <= io_input_payload_wr;
  io_outputs_0_payload_uncached <= io_input_payload_uncached;
  io_outputs_0_payload_address <= io_input_payload_address;
  io_outputs_0_payload_data <= io_input_payload_data;
  io_outputs_0_payload_mask <= io_input_payload_mask;
  io_outputs_0_payload_size <= io_input_payload_size;
  io_outputs_0_payload_last <= io_input_payload_last;
  io_outputs_0_fire <= (io_outputs_0_valid_read_buffer and io_outputs_0_ready);
  io_outputs_1_valid_read_buffer <= (io_input_valid and zz_io_outputs_1_valid);
  io_outputs_1_payload_wr <= io_input_payload_wr;
  io_outputs_1_payload_uncached <= io_input_payload_uncached;
  io_outputs_1_payload_address <= io_input_payload_address;
  io_outputs_1_payload_data <= io_input_payload_data;
  io_outputs_1_payload_mask <= io_input_payload_mask;
  io_outputs_1_payload_size <= io_input_payload_size;
  io_outputs_1_payload_last <= io_input_payload_last;
  io_outputs_1_fire <= (io_outputs_1_valid_read_buffer and io_outputs_1_ready);
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      zz_io_outputs_0_valid <= pkg_toStdLogic(true);
      zz_io_outputs_1_valid <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      if io_outputs_0_fire = '1' then
        zz_io_outputs_0_valid <= pkg_toStdLogic(false);
      end if;
      if io_outputs_1_fire = '1' then
        zz_io_outputs_1_valid <= pkg_toStdLogic(false);
      end if;
      if io_input_ready_read_buffer = '1' then
        zz_io_outputs_0_valid <= pkg_toStdLogic(true);
        zz_io_outputs_1_valid <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity JtagBridgeNoTap is
  port(
    io_ctrl_tdi : in std_logic;
    io_ctrl_enable : in std_logic;
    io_ctrl_capture : in std_logic;
    io_ctrl_shift : in std_logic;
    io_ctrl_update : in std_logic;
    io_ctrl_reset : in std_logic;
    io_ctrl_tdo : out std_logic;
    io_remote_cmd_valid : out std_logic;
    io_remote_cmd_ready : in std_logic;
    io_remote_cmd_payload_last : out std_logic;
    io_remote_cmd_payload_fragment : out std_logic_vector(0 downto 0);
    io_remote_rsp_valid : in std_logic;
    io_remote_rsp_ready : out std_logic;
    io_remote_rsp_payload_error : in std_logic;
    io_remote_rsp_payload_data : in std_logic_vector(31 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_systemReset : in std_logic;
    TCK : in std_logic
  );
end JtagBridgeNoTap;

architecture arch of JtagBridgeNoTap is
  signal io_remote_cmd_valid_read_buffer : std_logic;
  signal io_remote_rsp_ready_read_buffer : std_logic;
  signal flowCCByToggle_1_io_output_valid : std_logic;
  signal flowCCByToggle_1_io_output_payload_last : std_logic;
  signal flowCCByToggle_1_io_output_payload_fragment : std_logic_vector(0 downto 0);
  attribute async_reg : string;

  signal system_cmd_valid : std_logic;
  signal system_cmd_payload_last : std_logic;
  signal system_cmd_payload_fragment : std_logic_vector(0 downto 0);
  signal system_rsp_valid : std_logic;
  attribute async_reg of system_rsp_valid : signal is "true";
  signal system_rsp_payload_error : std_logic;
  attribute async_reg of system_rsp_payload_error : signal is "true";
  signal system_rsp_payload_data : std_logic_vector(31 downto 0);
  attribute async_reg of system_rsp_payload_data : signal is "true";
  signal io_remote_rsp_fire : std_logic;
  signal jtag_wrapper_ctrl_tdi : std_logic;
  signal jtag_wrapper_ctrl_enable : std_logic;
  signal jtag_wrapper_ctrl_capture : std_logic;
  signal jtag_wrapper_ctrl_shift : std_logic;
  signal jtag_wrapper_ctrl_update : std_logic;
  signal jtag_wrapper_ctrl_reset : std_logic;
  signal jtag_wrapper_ctrl_tdo : std_logic;
  signal jtag_wrapper_header : std_logic_vector(1 downto 0);
  signal jtag_wrapper_headerNext : std_logic_vector(1 downto 0);
  signal jtag_wrapper_counter : unsigned(0 downto 0);
  signal jtag_wrapper_done : std_logic;
  signal jtag_wrapper_sendCapture : std_logic;
  signal jtag_wrapper_sendShift : std_logic;
  signal jtag_wrapper_sendUpdate : std_logic;
  signal when_JtagTapInstructions_l185 : std_logic;
  signal when_JtagTapInstructions_l188 : std_logic;
  signal jtag_writeArea_ctrl_tdi : std_logic;
  signal jtag_writeArea_ctrl_enable : std_logic;
  signal jtag_writeArea_ctrl_capture : std_logic;
  signal jtag_writeArea_ctrl_shift : std_logic;
  signal jtag_writeArea_ctrl_update : std_logic;
  signal jtag_writeArea_ctrl_reset : std_logic;
  signal jtag_writeArea_ctrl_tdo : std_logic;
  signal jtag_writeArea_source_valid : std_logic;
  signal jtag_writeArea_source_payload_last : std_logic;
  signal jtag_writeArea_source_payload_fragment : std_logic_vector(0 downto 0);
  signal jtag_writeArea_valid : std_logic;
  signal jtag_writeArea_data : std_logic;
  signal when_JtagTapInstructions_l211 : std_logic;
  signal jtag_readArea_ctrl_tdi : std_logic;
  signal jtag_readArea_ctrl_enable : std_logic;
  signal jtag_readArea_ctrl_capture : std_logic;
  signal jtag_readArea_ctrl_shift : std_logic;
  signal jtag_readArea_ctrl_update : std_logic;
  signal jtag_readArea_ctrl_reset : std_logic;
  signal jtag_readArea_ctrl_tdo : std_logic;
  signal jtag_readArea_full_shifter : std_logic_vector(33 downto 0);
  signal when_JtagTapInstructions_l211_1 : std_logic;
begin
  io_remote_cmd_valid <= io_remote_cmd_valid_read_buffer;
  io_remote_rsp_ready <= io_remote_rsp_ready_read_buffer;
  flowCCByToggle_1 : entity work.FlowCCByToggle
    port map ( 
      io_input_valid => jtag_writeArea_source_valid,
      io_input_payload_last => jtag_writeArea_source_payload_last,
      io_input_payload_fragment => jtag_writeArea_source_payload_fragment,
      io_output_valid => flowCCByToggle_1_io_output_valid,
      io_output_payload_last => flowCCByToggle_1_io_output_payload_last,
      io_output_payload_fragment => flowCCByToggle_1_io_output_payload_fragment,
      TCK => TCK,
      io_mainClk => io_mainClk,
      resetCtrl_systemReset => resetCtrl_systemReset 
    );
  io_remote_cmd_valid_read_buffer <= system_cmd_valid;
  io_remote_cmd_payload_last <= system_cmd_payload_last;
  io_remote_cmd_payload_fragment <= system_cmd_payload_fragment;
  io_remote_rsp_fire <= (io_remote_rsp_valid and io_remote_rsp_ready_read_buffer);
  io_remote_rsp_ready_read_buffer <= pkg_toStdLogic(true);
  jtag_wrapper_headerNext <= pkg_shiftRight(pkg_cat(pkg_toStdLogicVector(jtag_wrapper_ctrl_tdi),jtag_wrapper_header),1);
  process(jtag_wrapper_ctrl_enable,jtag_wrapper_ctrl_shift,when_JtagTapInstructions_l185,when_JtagTapInstructions_l188)
  begin
    jtag_wrapper_sendCapture <= pkg_toStdLogic(false);
    if jtag_wrapper_ctrl_enable = '1' then
      if jtag_wrapper_ctrl_shift = '1' then
        if when_JtagTapInstructions_l185 = '1' then
          if when_JtagTapInstructions_l188 = '1' then
            jtag_wrapper_sendCapture <= pkg_toStdLogic(true);
          end if;
        end if;
      end if;
    end if;
  end process;

  process(jtag_wrapper_ctrl_enable,jtag_wrapper_ctrl_shift,when_JtagTapInstructions_l185)
  begin
    jtag_wrapper_sendShift <= pkg_toStdLogic(false);
    if jtag_wrapper_ctrl_enable = '1' then
      if jtag_wrapper_ctrl_shift = '1' then
        if when_JtagTapInstructions_l185 = '0' then
          jtag_wrapper_sendShift <= pkg_toStdLogic(true);
        end if;
      end if;
    end if;
  end process;

  process(jtag_wrapper_ctrl_enable,jtag_wrapper_ctrl_update)
  begin
    jtag_wrapper_sendUpdate <= pkg_toStdLogic(false);
    if jtag_wrapper_ctrl_enable = '1' then
      if jtag_wrapper_ctrl_update = '1' then
        jtag_wrapper_sendUpdate <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  when_JtagTapInstructions_l185 <= (not jtag_wrapper_done);
  when_JtagTapInstructions_l188 <= pkg_toStdLogic(jtag_wrapper_counter = pkg_unsigned("1"));
  process(when_JtagTapInstructions_l211,jtag_writeArea_ctrl_tdo,when_JtagTapInstructions_l211_1,jtag_readArea_ctrl_tdo)
  begin
    jtag_wrapper_ctrl_tdo <= pkg_toStdLogic(false);
    if when_JtagTapInstructions_l211 = '1' then
      jtag_wrapper_ctrl_tdo <= jtag_writeArea_ctrl_tdo;
    end if;
    if when_JtagTapInstructions_l211_1 = '1' then
      jtag_wrapper_ctrl_tdo <= jtag_readArea_ctrl_tdo;
    end if;
  end process;

  jtag_wrapper_ctrl_tdi <= io_ctrl_tdi;
  jtag_wrapper_ctrl_enable <= io_ctrl_enable;
  jtag_wrapper_ctrl_capture <= io_ctrl_capture;
  jtag_wrapper_ctrl_shift <= io_ctrl_shift;
  jtag_wrapper_ctrl_update <= io_ctrl_update;
  jtag_wrapper_ctrl_reset <= io_ctrl_reset;
  io_ctrl_tdo <= jtag_wrapper_ctrl_tdo;
  jtag_writeArea_source_valid <= jtag_writeArea_valid;
  jtag_writeArea_source_payload_last <= (not (jtag_writeArea_ctrl_enable and jtag_writeArea_ctrl_shift));
  jtag_writeArea_source_payload_fragment(0) <= jtag_writeArea_data;
  system_cmd_valid <= flowCCByToggle_1_io_output_valid;
  system_cmd_payload_last <= flowCCByToggle_1_io_output_payload_last;
  system_cmd_payload_fragment <= flowCCByToggle_1_io_output_payload_fragment;
  jtag_writeArea_ctrl_tdo <= pkg_toStdLogic(false);
  when_JtagTapInstructions_l211 <= pkg_toStdLogic(jtag_wrapper_header = pkg_stdLogicVector("00"));
  jtag_writeArea_ctrl_tdi <= jtag_wrapper_ctrl_tdi;
  jtag_writeArea_ctrl_enable <= pkg_toStdLogic(true);
  jtag_writeArea_ctrl_capture <= (pkg_toStdLogic(jtag_wrapper_headerNext = pkg_stdLogicVector("00")) and jtag_wrapper_sendCapture);
  jtag_writeArea_ctrl_shift <= (when_JtagTapInstructions_l211 and jtag_wrapper_sendShift);
  jtag_writeArea_ctrl_update <= (when_JtagTapInstructions_l211 and jtag_wrapper_sendUpdate);
  jtag_writeArea_ctrl_reset <= jtag_wrapper_ctrl_reset;
  jtag_readArea_ctrl_tdo <= pkg_extract(jtag_readArea_full_shifter,0);
  when_JtagTapInstructions_l211_1 <= pkg_toStdLogic(jtag_wrapper_header = pkg_stdLogicVector("01"));
  jtag_readArea_ctrl_tdi <= jtag_wrapper_ctrl_tdi;
  jtag_readArea_ctrl_enable <= pkg_toStdLogic(true);
  jtag_readArea_ctrl_capture <= (pkg_toStdLogic(jtag_wrapper_headerNext = pkg_stdLogicVector("01")) and jtag_wrapper_sendCapture);
  jtag_readArea_ctrl_shift <= (when_JtagTapInstructions_l211_1 and jtag_wrapper_sendShift);
  jtag_readArea_ctrl_update <= (when_JtagTapInstructions_l211_1 and jtag_wrapper_sendUpdate);
  jtag_readArea_ctrl_reset <= jtag_wrapper_ctrl_reset;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_remote_cmd_valid_read_buffer = '1' then
        system_rsp_valid <= pkg_toStdLogic(false);
      end if;
      if io_remote_rsp_fire = '1' then
        system_rsp_valid <= pkg_toStdLogic(true);
        system_rsp_payload_error <= io_remote_rsp_payload_error;
        system_rsp_payload_data <= io_remote_rsp_payload_data;
      end if;
    end if;
  end process;

  process(TCK)
  begin
    if rising_edge(TCK) then
      if jtag_wrapper_ctrl_enable = '1' then
        if jtag_wrapper_ctrl_capture = '1' then
          jtag_wrapper_done <= pkg_toStdLogic(false);
          jtag_wrapper_counter <= pkg_unsigned("0");
        end if;
        if jtag_wrapper_ctrl_shift = '1' then
          if when_JtagTapInstructions_l185 = '1' then
            jtag_wrapper_counter <= (jtag_wrapper_counter + pkg_unsigned("1"));
            jtag_wrapper_header <= jtag_wrapper_headerNext;
            if when_JtagTapInstructions_l188 = '1' then
              jtag_wrapper_done <= pkg_toStdLogic(true);
            end if;
          end if;
        end if;
      end if;
      jtag_writeArea_valid <= (jtag_writeArea_ctrl_enable and jtag_writeArea_ctrl_shift);
      jtag_writeArea_data <= jtag_writeArea_ctrl_tdi;
      if jtag_readArea_ctrl_enable = '1' then
        if jtag_readArea_ctrl_capture = '1' then
          jtag_readArea_full_shifter <= pkg_cat(pkg_cat(system_rsp_payload_data,pkg_toStdLogicVector(system_rsp_payload_error)),pkg_toStdLogicVector(system_rsp_valid));
        end if;
        if jtag_readArea_ctrl_shift = '1' then
          jtag_readArea_full_shifter <= pkg_shiftRight(pkg_cat(pkg_toStdLogicVector(jtag_readArea_ctrl_tdi),jtag_readArea_full_shifter),1);
        end if;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity SystemDebugger is
  port(
    io_remote_cmd_valid : in std_logic;
    io_remote_cmd_ready : out std_logic;
    io_remote_cmd_payload_last : in std_logic;
    io_remote_cmd_payload_fragment : in std_logic_vector(0 downto 0);
    io_remote_rsp_valid : out std_logic;
    io_remote_rsp_ready : in std_logic;
    io_remote_rsp_payload_error : out std_logic;
    io_remote_rsp_payload_data : out std_logic_vector(31 downto 0);
    io_mem_cmd_valid : out std_logic;
    io_mem_cmd_ready : in std_logic;
    io_mem_cmd_payload_address : out unsigned(31 downto 0);
    io_mem_cmd_payload_data : out std_logic_vector(31 downto 0);
    io_mem_cmd_payload_wr : out std_logic;
    io_mem_cmd_payload_size : out unsigned(1 downto 0);
    io_mem_rsp_valid : in std_logic;
    io_mem_rsp_payload : in std_logic_vector(31 downto 0);
    io_mainClk : in std_logic;
    resetCtrl_systemReset : in std_logic
  );
end SystemDebugger;

architecture arch of SystemDebugger is
  signal io_mem_cmd_valid_read_buffer : std_logic;

  signal dispatcher_dataShifter : std_logic_vector(66 downto 0);
  signal dispatcher_dataLoaded : std_logic;
  signal dispatcher_headerShifter : std_logic_vector(7 downto 0);
  signal dispatcher_header : std_logic_vector(7 downto 0);
  signal dispatcher_headerLoaded : std_logic;
  signal dispatcher_counter : unsigned(2 downto 0);
  signal when_Fragment_l346 : std_logic;
  signal when_Fragment_l349 : std_logic;
  signal zz_io_mem_cmd_payload_address : std_logic_vector(66 downto 0);
  signal io_mem_cmd_isStall : std_logic;
  signal when_Fragment_l372 : std_logic;
begin
  io_mem_cmd_valid <= io_mem_cmd_valid_read_buffer;
  dispatcher_header <= pkg_extract(dispatcher_headerShifter,7,0);
  when_Fragment_l346 <= pkg_toStdLogic(dispatcher_headerLoaded = pkg_toStdLogic(false));
  when_Fragment_l349 <= pkg_toStdLogic(dispatcher_counter = pkg_unsigned("111"));
  io_remote_cmd_ready <= (not dispatcher_dataLoaded);
  zz_io_mem_cmd_payload_address <= pkg_extract(dispatcher_dataShifter,66,0);
  io_mem_cmd_payload_address <= unsigned(pkg_extract(zz_io_mem_cmd_payload_address,31,0));
  io_mem_cmd_payload_data <= pkg_extract(zz_io_mem_cmd_payload_address,63,32);
  io_mem_cmd_payload_wr <= pkg_extract(zz_io_mem_cmd_payload_address,64);
  io_mem_cmd_payload_size <= unsigned(pkg_extract(zz_io_mem_cmd_payload_address,66,65));
  io_mem_cmd_valid_read_buffer <= (dispatcher_dataLoaded and pkg_toStdLogic(dispatcher_header = pkg_stdLogicVector("00000000")));
  io_mem_cmd_isStall <= (io_mem_cmd_valid_read_buffer and (not io_mem_cmd_ready));
  when_Fragment_l372 <= ((dispatcher_headerLoaded and dispatcher_dataLoaded) and (not io_mem_cmd_isStall));
  io_remote_rsp_valid <= io_mem_rsp_valid;
  io_remote_rsp_payload_error <= pkg_toStdLogic(false);
  io_remote_rsp_payload_data <= io_mem_rsp_payload;
  process(io_mainClk, resetCtrl_systemReset)
  begin
    if resetCtrl_systemReset = '1' then
      dispatcher_dataLoaded <= pkg_toStdLogic(false);
      dispatcher_headerLoaded <= pkg_toStdLogic(false);
      dispatcher_counter <= pkg_unsigned("000");
    elsif rising_edge(io_mainClk) then
      if io_remote_cmd_valid = '1' then
        if when_Fragment_l346 = '1' then
          dispatcher_counter <= (dispatcher_counter + pkg_unsigned("001"));
          if when_Fragment_l349 = '1' then
            dispatcher_headerLoaded <= pkg_toStdLogic(true);
          end if;
        end if;
        if io_remote_cmd_payload_last = '1' then
          dispatcher_headerLoaded <= pkg_toStdLogic(true);
          dispatcher_dataLoaded <= pkg_toStdLogic(true);
          dispatcher_counter <= pkg_unsigned("000");
        end if;
      end if;
      if when_Fragment_l372 = '1' then
        dispatcher_headerLoaded <= pkg_toStdLogic(false);
        dispatcher_dataLoaded <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if io_remote_cmd_valid = '1' then
        if when_Fragment_l346 = '1' then
          dispatcher_headerShifter <= pkg_shiftRight(pkg_cat(io_remote_cmd_payload_fragment,dispatcher_headerShifter),1);
        else
          dispatcher_dataShifter <= pkg_shiftRight(pkg_cat(io_remote_cmd_payload_fragment,dispatcher_dataShifter),1);
        end if;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4ReadOnlyDecoder is
  port(
    io_input_ar_valid : in std_logic;
    io_input_ar_ready : out std_logic;
    io_input_ar_payload_addr : in unsigned(31 downto 0);
    io_input_ar_payload_len : in unsigned(7 downto 0);
    io_input_ar_payload_burst : in std_logic_vector(1 downto 0);
    io_input_ar_payload_cache : in std_logic_vector(3 downto 0);
    io_input_ar_payload_prot : in std_logic_vector(2 downto 0);
    io_input_r_valid : out std_logic;
    io_input_r_ready : in std_logic;
    io_input_r_payload_data : out std_logic_vector(31 downto 0);
    io_input_r_payload_resp : out std_logic_vector(1 downto 0);
    io_input_r_payload_last : out std_logic;
    io_outputs_0_ar_valid : out std_logic;
    io_outputs_0_ar_ready : in std_logic;
    io_outputs_0_ar_payload_addr : out unsigned(31 downto 0);
    io_outputs_0_ar_payload_len : out unsigned(7 downto 0);
    io_outputs_0_ar_payload_burst : out std_logic_vector(1 downto 0);
    io_outputs_0_ar_payload_cache : out std_logic_vector(3 downto 0);
    io_outputs_0_ar_payload_prot : out std_logic_vector(2 downto 0);
    io_outputs_0_r_valid : in std_logic;
    io_outputs_0_r_ready : out std_logic;
    io_outputs_0_r_payload_data : in std_logic_vector(31 downto 0);
    io_outputs_0_r_payload_resp : in std_logic_vector(1 downto 0);
    io_outputs_0_r_payload_last : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4ReadOnlyDecoder;

architecture arch of Axi4ReadOnlyDecoder is
  signal errorSlave_io_axi_ar_valid : std_logic;
  signal io_input_ar_ready_read_buffer : std_logic;
  signal io_input_r_valid_read_buffer : std_logic;
  signal io_input_r_payload_last_read_buffer : std_logic;
  signal errorSlave_io_axi_ar_ready : std_logic;
  signal errorSlave_io_axi_r_valid : std_logic;
  signal errorSlave_io_axi_r_payload_data : std_logic_vector(31 downto 0);
  signal errorSlave_io_axi_r_payload_resp : std_logic_vector(1 downto 0);
  signal errorSlave_io_axi_r_payload_last : std_logic;

  signal io_input_ar_fire : std_logic;
  signal io_input_r_fire : std_logic;
  signal when_Utils_l597 : std_logic;
  signal pendingCmdCounter_incrementIt : std_logic;
  signal pendingCmdCounter_decrementIt : std_logic;
  signal pendingCmdCounter_valueNext : unsigned(2 downto 0);
  signal pendingCmdCounter_value : unsigned(2 downto 0);
  signal pendingCmdCounter_willOverflowIfInc : std_logic;
  signal pendingCmdCounter_willOverflow : std_logic;
  signal pendingCmdCounter_finalIncrement : unsigned(2 downto 0);
  signal when_Utils_l622 : std_logic;
  signal when_Utils_l624 : std_logic;
  signal decodedCmdSels : std_logic_vector(0 downto 0);
  signal decodedCmdError : std_logic;
  signal pendingSels : std_logic_vector(0 downto 0);
  signal pendingError : std_logic;
  signal allowCmd : std_logic;
begin
  io_input_ar_ready <= io_input_ar_ready_read_buffer;
  io_input_r_valid <= io_input_r_valid_read_buffer;
  io_input_r_payload_last <= io_input_r_payload_last_read_buffer;
  errorSlave : entity work.Axi4ReadOnlyErrorSlave
    port map ( 
      io_axi_ar_valid => errorSlave_io_axi_ar_valid,
      io_axi_ar_ready => errorSlave_io_axi_ar_ready,
      io_axi_ar_payload_addr => io_input_ar_payload_addr,
      io_axi_ar_payload_len => io_input_ar_payload_len,
      io_axi_ar_payload_burst => io_input_ar_payload_burst,
      io_axi_ar_payload_cache => io_input_ar_payload_cache,
      io_axi_ar_payload_prot => io_input_ar_payload_prot,
      io_axi_r_valid => errorSlave_io_axi_r_valid,
      io_axi_r_ready => io_input_r_ready,
      io_axi_r_payload_data => errorSlave_io_axi_r_payload_data,
      io_axi_r_payload_resp => errorSlave_io_axi_r_payload_resp,
      io_axi_r_payload_last => errorSlave_io_axi_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  io_input_ar_fire <= (io_input_ar_valid and io_input_ar_ready_read_buffer);
  io_input_r_fire <= (io_input_r_valid_read_buffer and io_input_r_ready);
  when_Utils_l597 <= (io_input_r_fire and io_input_r_payload_last_read_buffer);
  process(io_input_ar_fire)
  begin
    pendingCmdCounter_incrementIt <= pkg_toStdLogic(false);
    if io_input_ar_fire = '1' then
      pendingCmdCounter_incrementIt <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_Utils_l597)
  begin
    pendingCmdCounter_decrementIt <= pkg_toStdLogic(false);
    if when_Utils_l597 = '1' then
      pendingCmdCounter_decrementIt <= pkg_toStdLogic(true);
    end if;
  end process;

  pendingCmdCounter_willOverflowIfInc <= (pkg_toStdLogic(pendingCmdCounter_value = pkg_unsigned("111")) and (not pendingCmdCounter_decrementIt));
  pendingCmdCounter_willOverflow <= (pendingCmdCounter_willOverflowIfInc and pendingCmdCounter_incrementIt);
  when_Utils_l622 <= (pendingCmdCounter_incrementIt and (not pendingCmdCounter_decrementIt));
  process(when_Utils_l622,when_Utils_l624)
  begin
    if when_Utils_l622 = '1' then
      pendingCmdCounter_finalIncrement <= pkg_unsigned("001");
    else
      if when_Utils_l624 = '1' then
        pendingCmdCounter_finalIncrement <= pkg_unsigned("111");
      else
        pendingCmdCounter_finalIncrement <= pkg_unsigned("000");
      end if;
    end if;
  end process;

  when_Utils_l624 <= ((not pendingCmdCounter_incrementIt) and pendingCmdCounter_decrementIt);
  pendingCmdCounter_valueNext <= (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  decodedCmdSels <= pkg_toStdLogicVector((pkg_toStdLogic((io_input_ar_payload_addr and pkg_not(pkg_unsigned("00000000000000000111111111111111"))) = pkg_unsigned("10000000000000000000000000000000")) and io_input_ar_valid));
  decodedCmdError <= pkg_toStdLogic(decodedCmdSels = pkg_stdLogicVector("0"));
  allowCmd <= (pkg_toStdLogic(pendingCmdCounter_value = pkg_unsigned("000")) or (pkg_toStdLogic(pendingCmdCounter_value /= pkg_unsigned("111")) and pkg_toStdLogic(pendingSels = decodedCmdSels)));
  io_input_ar_ready_read_buffer <= ((pkg_toStdLogic((decodedCmdSels and pkg_toStdLogicVector(io_outputs_0_ar_ready)) /= pkg_stdLogicVector("0")) or (decodedCmdError and errorSlave_io_axi_ar_ready)) and allowCmd);
  errorSlave_io_axi_ar_valid <= ((io_input_ar_valid and decodedCmdError) and allowCmd);
  io_outputs_0_ar_valid <= ((io_input_ar_valid and pkg_extract(decodedCmdSels,0)) and allowCmd);
  io_outputs_0_ar_payload_addr <= io_input_ar_payload_addr;
  io_outputs_0_ar_payload_len <= io_input_ar_payload_len;
  io_outputs_0_ar_payload_burst <= io_input_ar_payload_burst;
  io_outputs_0_ar_payload_cache <= io_input_ar_payload_cache;
  io_outputs_0_ar_payload_prot <= io_input_ar_payload_prot;
  process(io_outputs_0_r_valid,errorSlave_io_axi_r_valid)
  begin
    io_input_r_valid_read_buffer <= pkg_toStdLogic(pkg_toStdLogicVector(io_outputs_0_r_valid) /= pkg_stdLogicVector("0"));
    if errorSlave_io_axi_r_valid = '1' then
      io_input_r_valid_read_buffer <= pkg_toStdLogic(true);
    end if;
  end process;

  io_input_r_payload_data <= io_outputs_0_r_payload_data;
  process(io_outputs_0_r_payload_resp,pendingError,errorSlave_io_axi_r_payload_resp)
  begin
    io_input_r_payload_resp <= io_outputs_0_r_payload_resp;
    if pendingError = '1' then
      io_input_r_payload_resp <= errorSlave_io_axi_r_payload_resp;
    end if;
  end process;

  process(io_outputs_0_r_payload_last,pendingError,errorSlave_io_axi_r_payload_last)
  begin
    io_input_r_payload_last_read_buffer <= io_outputs_0_r_payload_last;
    if pendingError = '1' then
      io_input_r_payload_last_read_buffer <= errorSlave_io_axi_r_payload_last;
    end if;
  end process;

  io_outputs_0_r_ready <= io_input_r_ready;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      pendingCmdCounter_value <= pkg_unsigned("000");
      pendingSels <= pkg_stdLogicVector("0");
      pendingError <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      if io_input_ar_ready_read_buffer = '1' then
        pendingSels <= decodedCmdSels;
      end if;
      if io_input_ar_ready_read_buffer = '1' then
        pendingError <= decodedCmdError;
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4SharedDecoder is
  port(
    io_input_arw_valid : in std_logic;
    io_input_arw_ready : out std_logic;
    io_input_arw_payload_addr : in unsigned(31 downto 0);
    io_input_arw_payload_len : in unsigned(7 downto 0);
    io_input_arw_payload_size : in unsigned(2 downto 0);
    io_input_arw_payload_cache : in std_logic_vector(3 downto 0);
    io_input_arw_payload_prot : in std_logic_vector(2 downto 0);
    io_input_arw_payload_write : in std_logic;
    io_input_w_valid : in std_logic;
    io_input_w_ready : out std_logic;
    io_input_w_payload_data : in std_logic_vector(31 downto 0);
    io_input_w_payload_strb : in std_logic_vector(3 downto 0);
    io_input_w_payload_last : in std_logic;
    io_input_b_valid : out std_logic;
    io_input_b_ready : in std_logic;
    io_input_b_payload_resp : out std_logic_vector(1 downto 0);
    io_input_r_valid : out std_logic;
    io_input_r_ready : in std_logic;
    io_input_r_payload_data : out std_logic_vector(31 downto 0);
    io_input_r_payload_resp : out std_logic_vector(1 downto 0);
    io_input_r_payload_last : out std_logic;
    io_sharedOutputs_0_arw_valid : out std_logic;
    io_sharedOutputs_0_arw_ready : in std_logic;
    io_sharedOutputs_0_arw_payload_addr : out unsigned(31 downto 0);
    io_sharedOutputs_0_arw_payload_len : out unsigned(7 downto 0);
    io_sharedOutputs_0_arw_payload_size : out unsigned(2 downto 0);
    io_sharedOutputs_0_arw_payload_cache : out std_logic_vector(3 downto 0);
    io_sharedOutputs_0_arw_payload_prot : out std_logic_vector(2 downto 0);
    io_sharedOutputs_0_arw_payload_write : out std_logic;
    io_sharedOutputs_0_w_valid : out std_logic;
    io_sharedOutputs_0_w_ready : in std_logic;
    io_sharedOutputs_0_w_payload_data : out std_logic_vector(31 downto 0);
    io_sharedOutputs_0_w_payload_strb : out std_logic_vector(3 downto 0);
    io_sharedOutputs_0_w_payload_last : out std_logic;
    io_sharedOutputs_0_b_valid : in std_logic;
    io_sharedOutputs_0_b_ready : out std_logic;
    io_sharedOutputs_0_b_payload_resp : in std_logic_vector(1 downto 0);
    io_sharedOutputs_0_r_valid : in std_logic;
    io_sharedOutputs_0_r_ready : out std_logic;
    io_sharedOutputs_0_r_payload_data : in std_logic_vector(31 downto 0);
    io_sharedOutputs_0_r_payload_resp : in std_logic_vector(1 downto 0);
    io_sharedOutputs_0_r_payload_last : in std_logic;
    io_sharedOutputs_1_arw_valid : out std_logic;
    io_sharedOutputs_1_arw_ready : in std_logic;
    io_sharedOutputs_1_arw_payload_addr : out unsigned(31 downto 0);
    io_sharedOutputs_1_arw_payload_len : out unsigned(7 downto 0);
    io_sharedOutputs_1_arw_payload_size : out unsigned(2 downto 0);
    io_sharedOutputs_1_arw_payload_cache : out std_logic_vector(3 downto 0);
    io_sharedOutputs_1_arw_payload_prot : out std_logic_vector(2 downto 0);
    io_sharedOutputs_1_arw_payload_write : out std_logic;
    io_sharedOutputs_1_w_valid : out std_logic;
    io_sharedOutputs_1_w_ready : in std_logic;
    io_sharedOutputs_1_w_payload_data : out std_logic_vector(31 downto 0);
    io_sharedOutputs_1_w_payload_strb : out std_logic_vector(3 downto 0);
    io_sharedOutputs_1_w_payload_last : out std_logic;
    io_sharedOutputs_1_b_valid : in std_logic;
    io_sharedOutputs_1_b_ready : out std_logic;
    io_sharedOutputs_1_b_payload_resp : in std_logic_vector(1 downto 0);
    io_sharedOutputs_1_r_valid : in std_logic;
    io_sharedOutputs_1_r_ready : out std_logic;
    io_sharedOutputs_1_r_payload_data : in std_logic_vector(31 downto 0);
    io_sharedOutputs_1_r_payload_resp : in std_logic_vector(1 downto 0);
    io_sharedOutputs_1_r_payload_last : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4SharedDecoder;

architecture arch of Axi4SharedDecoder is
  signal errorSlave_io_axi_arw_valid : std_logic;
  signal errorSlave_io_axi_w_valid : std_logic;
  signal io_input_arw_ready_read_buffer : std_logic;
  signal io_input_b_valid_read_buffer : std_logic;
  signal io_input_r_valid_read_buffer : std_logic;
  signal io_input_r_payload_last_read_buffer : std_logic;
  signal io_input_w_ready_read_buffer : std_logic;
  signal errorSlave_io_axi_arw_ready : std_logic;
  signal errorSlave_io_axi_w_ready : std_logic;
  signal errorSlave_io_axi_b_valid : std_logic;
  signal errorSlave_io_axi_b_payload_resp : std_logic_vector(1 downto 0);
  signal errorSlave_io_axi_r_valid : std_logic;
  signal errorSlave_io_axi_r_payload_data : std_logic_vector(31 downto 0);
  signal errorSlave_io_axi_r_payload_resp : std_logic_vector(1 downto 0);
  signal errorSlave_io_axi_r_payload_last : std_logic;
  signal zz_io_input_b_payload_resp : std_logic_vector(1 downto 0);
  signal zz_io_input_r_payload_data : std_logic_vector(31 downto 0);
  signal zz_io_input_r_payload_resp : std_logic_vector(1 downto 0);
  signal zz_io_input_r_payload_last : std_logic;

  signal zz_pendingCmdCounter : unsigned(2 downto 0);
  signal zz_pendingCmdCounter_1 : unsigned(2 downto 0);
  signal zz_pendingCmdCounter_2 : unsigned(2 downto 0);
  signal cmdAllowedStart : std_logic;
  signal io_input_arw_fire : std_logic;
  signal io_input_b_fire : std_logic;
  signal io_input_r_fire : std_logic;
  signal when_Utils_l648 : std_logic;
  signal pendingCmdCounter : unsigned(2 downto 0);
  signal zz_pendingCmdCounter_3 : unsigned(2 downto 0);
  signal when_Utils_l594 : std_logic;
  signal io_input_w_fire : std_logic;
  signal when_Utils_l597 : std_logic;
  signal pendingDataCounter_incrementIt : std_logic;
  signal pendingDataCounter_decrementIt : std_logic;
  signal pendingDataCounter_valueNext : unsigned(2 downto 0);
  signal pendingDataCounter_value : unsigned(2 downto 0);
  signal pendingDataCounter_willOverflowIfInc : std_logic;
  signal pendingDataCounter_willOverflow : std_logic;
  signal pendingDataCounter_finalIncrement : unsigned(2 downto 0);
  signal when_Utils_l622 : std_logic;
  signal when_Utils_l624 : std_logic;
  signal decodedCmdSels : std_logic_vector(1 downto 0);
  signal decodedCmdError : std_logic;
  signal pendingSels : std_logic_vector(1 downto 0);
  signal pendingError : std_logic;
  signal allowCmd : std_logic;
  signal allowData : std_logic;
  signal zz_cmdAllowedStart : std_logic;
  signal zz_io_sharedOutputs_0_arw_valid : std_logic_vector(1 downto 0);
  signal zz_io_sharedOutputs_0_w_valid : std_logic_vector(1 downto 0);
  signal zz_writeRspIndex : std_logic;
  signal writeRspIndex : unsigned(0 downto 0);
  signal zz_readRspIndex : std_logic;
  signal readRspIndex : unsigned(0 downto 0);
begin
  io_input_arw_ready <= io_input_arw_ready_read_buffer;
  io_input_b_valid <= io_input_b_valid_read_buffer;
  io_input_r_valid <= io_input_r_valid_read_buffer;
  io_input_r_payload_last <= io_input_r_payload_last_read_buffer;
  io_input_w_ready <= io_input_w_ready_read_buffer;
  errorSlave : entity work.Axi4SharedErrorSlave
    port map ( 
      io_axi_arw_valid => errorSlave_io_axi_arw_valid,
      io_axi_arw_ready => errorSlave_io_axi_arw_ready,
      io_axi_arw_payload_addr => io_input_arw_payload_addr,
      io_axi_arw_payload_len => io_input_arw_payload_len,
      io_axi_arw_payload_size => io_input_arw_payload_size,
      io_axi_arw_payload_cache => io_input_arw_payload_cache,
      io_axi_arw_payload_prot => io_input_arw_payload_prot,
      io_axi_arw_payload_write => io_input_arw_payload_write,
      io_axi_w_valid => errorSlave_io_axi_w_valid,
      io_axi_w_ready => errorSlave_io_axi_w_ready,
      io_axi_w_payload_data => io_input_w_payload_data,
      io_axi_w_payload_strb => io_input_w_payload_strb,
      io_axi_w_payload_last => io_input_w_payload_last,
      io_axi_b_valid => errorSlave_io_axi_b_valid,
      io_axi_b_ready => io_input_b_ready,
      io_axi_b_payload_resp => errorSlave_io_axi_b_payload_resp,
      io_axi_r_valid => errorSlave_io_axi_r_valid,
      io_axi_r_ready => io_input_r_ready,
      io_axi_r_payload_data => errorSlave_io_axi_r_payload_data,
      io_axi_r_payload_resp => errorSlave_io_axi_r_payload_resp,
      io_axi_r_payload_last => errorSlave_io_axi_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  process(writeRspIndex,io_sharedOutputs_0_b_payload_resp,io_sharedOutputs_1_b_payload_resp)
  begin
    case writeRspIndex is
      when "0" =>
        zz_io_input_b_payload_resp <= io_sharedOutputs_0_b_payload_resp;
      when others =>
        zz_io_input_b_payload_resp <= io_sharedOutputs_1_b_payload_resp;
    end case;
  end process;

  process(readRspIndex,io_sharedOutputs_0_r_payload_data,io_sharedOutputs_0_r_payload_resp,io_sharedOutputs_0_r_payload_last,io_sharedOutputs_1_r_payload_data,io_sharedOutputs_1_r_payload_resp,io_sharedOutputs_1_r_payload_last)
  begin
    case readRspIndex is
      when "0" =>
        zz_io_input_r_payload_data <= io_sharedOutputs_0_r_payload_data;
        zz_io_input_r_payload_resp <= io_sharedOutputs_0_r_payload_resp;
        zz_io_input_r_payload_last <= io_sharedOutputs_0_r_payload_last;
      when others =>
        zz_io_input_r_payload_data <= io_sharedOutputs_1_r_payload_data;
        zz_io_input_r_payload_resp <= io_sharedOutputs_1_r_payload_resp;
        zz_io_input_r_payload_last <= io_sharedOutputs_1_r_payload_last;
    end case;
  end process;

  process(zz_pendingCmdCounter_1,when_Utils_l648)
  begin
    zz_pendingCmdCounter <= zz_pendingCmdCounter_1;
    if when_Utils_l648 = '1' then
      zz_pendingCmdCounter <= (zz_pendingCmdCounter_1 - pkg_unsigned("001"));
    end if;
  end process;

  process(zz_pendingCmdCounter_2,io_input_b_fire)
  begin
    zz_pendingCmdCounter_1 <= zz_pendingCmdCounter_2;
    if io_input_b_fire = '1' then
      zz_pendingCmdCounter_1 <= (zz_pendingCmdCounter_2 - pkg_unsigned("001"));
    end if;
  end process;

  process(zz_pendingCmdCounter_3,io_input_arw_fire)
  begin
    zz_pendingCmdCounter_2 <= zz_pendingCmdCounter_3;
    if io_input_arw_fire = '1' then
      zz_pendingCmdCounter_2 <= (zz_pendingCmdCounter_3 + pkg_unsigned("001"));
    end if;
  end process;

  io_input_arw_fire <= (io_input_arw_valid and io_input_arw_ready_read_buffer);
  io_input_b_fire <= (io_input_b_valid_read_buffer and io_input_b_ready);
  io_input_r_fire <= (io_input_r_valid_read_buffer and io_input_r_ready);
  when_Utils_l648 <= (io_input_r_fire and io_input_r_payload_last_read_buffer);
  zz_pendingCmdCounter_3 <= pendingCmdCounter;
  when_Utils_l594 <= (cmdAllowedStart and io_input_arw_payload_write);
  io_input_w_fire <= (io_input_w_valid and io_input_w_ready_read_buffer);
  when_Utils_l597 <= (io_input_w_fire and io_input_w_payload_last);
  process(when_Utils_l594)
  begin
    pendingDataCounter_incrementIt <= pkg_toStdLogic(false);
    if when_Utils_l594 = '1' then
      pendingDataCounter_incrementIt <= pkg_toStdLogic(true);
    end if;
  end process;

  process(when_Utils_l597)
  begin
    pendingDataCounter_decrementIt <= pkg_toStdLogic(false);
    if when_Utils_l597 = '1' then
      pendingDataCounter_decrementIt <= pkg_toStdLogic(true);
    end if;
  end process;

  pendingDataCounter_willOverflowIfInc <= (pkg_toStdLogic(pendingDataCounter_value = pkg_unsigned("111")) and (not pendingDataCounter_decrementIt));
  pendingDataCounter_willOverflow <= (pendingDataCounter_willOverflowIfInc and pendingDataCounter_incrementIt);
  when_Utils_l622 <= (pendingDataCounter_incrementIt and (not pendingDataCounter_decrementIt));
  process(when_Utils_l622,when_Utils_l624)
  begin
    if when_Utils_l622 = '1' then
      pendingDataCounter_finalIncrement <= pkg_unsigned("001");
    else
      if when_Utils_l624 = '1' then
        pendingDataCounter_finalIncrement <= pkg_unsigned("111");
      else
        pendingDataCounter_finalIncrement <= pkg_unsigned("000");
      end if;
    end if;
  end process;

  when_Utils_l624 <= ((not pendingDataCounter_incrementIt) and pendingDataCounter_decrementIt);
  pendingDataCounter_valueNext <= (pendingDataCounter_value + pendingDataCounter_finalIncrement);
  decodedCmdSels <= pkg_cat(pkg_toStdLogicVector(pkg_toStdLogic((io_input_arw_payload_addr and pkg_not(pkg_unsigned("00000000000011111111111111111111"))) = pkg_unsigned("11110000000000000000000000000000"))),pkg_toStdLogicVector(pkg_toStdLogic((io_input_arw_payload_addr and pkg_not(pkg_unsigned("00000000000000000111111111111111"))) = pkg_unsigned("10000000000000000000000000000000"))));
  decodedCmdError <= pkg_toStdLogic(decodedCmdSels = pkg_stdLogicVector("00"));
  allowCmd <= (pkg_toStdLogic(pendingCmdCounter = pkg_unsigned("000")) or (pkg_toStdLogic(pendingCmdCounter /= pkg_unsigned("111")) and pkg_toStdLogic(pendingSels = decodedCmdSels)));
  allowData <= pkg_toStdLogic(pendingDataCounter_value /= pkg_unsigned("000"));
  cmdAllowedStart <= ((io_input_arw_valid and allowCmd) and zz_cmdAllowedStart);
  io_input_arw_ready_read_buffer <= ((pkg_toStdLogic((decodedCmdSels and pkg_cat(pkg_toStdLogicVector(io_sharedOutputs_1_arw_ready),pkg_toStdLogicVector(io_sharedOutputs_0_arw_ready))) /= pkg_stdLogicVector("00")) or (decodedCmdError and errorSlave_io_axi_arw_ready)) and allowCmd);
  errorSlave_io_axi_arw_valid <= ((io_input_arw_valid and decodedCmdError) and allowCmd);
  zz_io_sharedOutputs_0_arw_valid <= pkg_extract(decodedCmdSels,1,0);
  io_sharedOutputs_0_arw_valid <= ((io_input_arw_valid and pkg_extract(zz_io_sharedOutputs_0_arw_valid,0)) and allowCmd);
  io_sharedOutputs_0_arw_payload_addr <= io_input_arw_payload_addr;
  io_sharedOutputs_0_arw_payload_len <= io_input_arw_payload_len;
  io_sharedOutputs_0_arw_payload_size <= io_input_arw_payload_size;
  io_sharedOutputs_0_arw_payload_cache <= io_input_arw_payload_cache;
  io_sharedOutputs_0_arw_payload_prot <= io_input_arw_payload_prot;
  io_sharedOutputs_0_arw_payload_write <= io_input_arw_payload_write;
  io_sharedOutputs_1_arw_valid <= ((io_input_arw_valid and pkg_extract(zz_io_sharedOutputs_0_arw_valid,1)) and allowCmd);
  io_sharedOutputs_1_arw_payload_addr <= io_input_arw_payload_addr;
  io_sharedOutputs_1_arw_payload_len <= io_input_arw_payload_len;
  io_sharedOutputs_1_arw_payload_size <= io_input_arw_payload_size;
  io_sharedOutputs_1_arw_payload_cache <= io_input_arw_payload_cache;
  io_sharedOutputs_1_arw_payload_prot <= io_input_arw_payload_prot;
  io_sharedOutputs_1_arw_payload_write <= io_input_arw_payload_write;
  io_input_w_ready_read_buffer <= ((pkg_toStdLogic((pkg_extract(pendingSels,1,0) and pkg_cat(pkg_toStdLogicVector(io_sharedOutputs_1_w_ready),pkg_toStdLogicVector(io_sharedOutputs_0_w_ready))) /= pkg_stdLogicVector("00")) or (pendingError and errorSlave_io_axi_w_ready)) and allowData);
  errorSlave_io_axi_w_valid <= ((io_input_w_valid and pendingError) and allowData);
  zz_io_sharedOutputs_0_w_valid <= pkg_extract(pendingSels,1,0);
  io_sharedOutputs_0_w_valid <= ((io_input_w_valid and pkg_extract(zz_io_sharedOutputs_0_w_valid,0)) and allowData);
  io_sharedOutputs_0_w_payload_data <= io_input_w_payload_data;
  io_sharedOutputs_0_w_payload_strb <= io_input_w_payload_strb;
  io_sharedOutputs_0_w_payload_last <= io_input_w_payload_last;
  io_sharedOutputs_1_w_valid <= ((io_input_w_valid and pkg_extract(zz_io_sharedOutputs_0_w_valid,1)) and allowData);
  io_sharedOutputs_1_w_payload_data <= io_input_w_payload_data;
  io_sharedOutputs_1_w_payload_strb <= io_input_w_payload_strb;
  io_sharedOutputs_1_w_payload_last <= io_input_w_payload_last;
  zz_writeRspIndex <= pkg_extract(pkg_extract(pendingSels,1,0),1);
  writeRspIndex <= unsigned(pkg_toStdLogicVector(zz_writeRspIndex));
  io_input_b_valid_read_buffer <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(io_sharedOutputs_1_b_valid),pkg_toStdLogicVector(io_sharedOutputs_0_b_valid)) /= pkg_stdLogicVector("00")) or errorSlave_io_axi_b_valid);
  process(zz_io_input_b_payload_resp,pendingError,errorSlave_io_axi_b_payload_resp)
  begin
    io_input_b_payload_resp <= zz_io_input_b_payload_resp;
    if pendingError = '1' then
      io_input_b_payload_resp <= errorSlave_io_axi_b_payload_resp;
    end if;
  end process;

  io_sharedOutputs_0_b_ready <= io_input_b_ready;
  io_sharedOutputs_1_b_ready <= io_input_b_ready;
  zz_readRspIndex <= pkg_extract(pkg_extract(pendingSels,1,0),1);
  readRspIndex <= unsigned(pkg_toStdLogicVector(zz_readRspIndex));
  io_input_r_valid_read_buffer <= (pkg_toStdLogic(pkg_cat(pkg_toStdLogicVector(io_sharedOutputs_1_r_valid),pkg_toStdLogicVector(io_sharedOutputs_0_r_valid)) /= pkg_stdLogicVector("00")) or errorSlave_io_axi_r_valid);
  io_input_r_payload_data <= zz_io_input_r_payload_data;
  process(zz_io_input_r_payload_resp,pendingError,errorSlave_io_axi_r_payload_resp)
  begin
    io_input_r_payload_resp <= zz_io_input_r_payload_resp;
    if pendingError = '1' then
      io_input_r_payload_resp <= errorSlave_io_axi_r_payload_resp;
    end if;
  end process;

  process(zz_io_input_r_payload_last,pendingError,errorSlave_io_axi_r_payload_last)
  begin
    io_input_r_payload_last_read_buffer <= zz_io_input_r_payload_last;
    if pendingError = '1' then
      io_input_r_payload_last_read_buffer <= errorSlave_io_axi_r_payload_last;
    end if;
  end process;

  io_sharedOutputs_0_r_ready <= io_input_r_ready;
  io_sharedOutputs_1_r_ready <= io_input_r_ready;
  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      pendingCmdCounter <= pkg_unsigned("000");
      pendingDataCounter_value <= pkg_unsigned("000");
      pendingSels <= pkg_stdLogicVector("00");
      pendingError <= pkg_toStdLogic(false);
      zz_cmdAllowedStart <= pkg_toStdLogic(true);
    elsif rising_edge(io_mainClk) then
      pendingCmdCounter <= zz_pendingCmdCounter;
      pendingDataCounter_value <= pendingDataCounter_valueNext;
      if cmdAllowedStart = '1' then
        pendingSels <= decodedCmdSels;
      end if;
      if cmdAllowedStart = '1' then
        pendingError <= decodedCmdError;
      end if;
      if cmdAllowedStart = '1' then
        zz_cmdAllowedStart <= pkg_toStdLogic(false);
      end if;
      if io_input_arw_ready_read_buffer = '1' then
        zz_cmdAllowedStart <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4SharedArbiter is
  port(
    io_readInputs_0_ar_valid : in std_logic;
    io_readInputs_0_ar_ready : out std_logic;
    io_readInputs_0_ar_payload_addr : in unsigned(14 downto 0);
    io_readInputs_0_ar_payload_id : in unsigned(2 downto 0);
    io_readInputs_0_ar_payload_len : in unsigned(7 downto 0);
    io_readInputs_0_ar_payload_size : in unsigned(2 downto 0);
    io_readInputs_0_ar_payload_burst : in std_logic_vector(1 downto 0);
    io_readInputs_0_r_valid : out std_logic;
    io_readInputs_0_r_ready : in std_logic;
    io_readInputs_0_r_payload_data : out std_logic_vector(31 downto 0);
    io_readInputs_0_r_payload_id : out unsigned(2 downto 0);
    io_readInputs_0_r_payload_resp : out std_logic_vector(1 downto 0);
    io_readInputs_0_r_payload_last : out std_logic;
    io_sharedInputs_0_arw_valid : in std_logic;
    io_sharedInputs_0_arw_ready : out std_logic;
    io_sharedInputs_0_arw_payload_addr : in unsigned(14 downto 0);
    io_sharedInputs_0_arw_payload_id : in unsigned(2 downto 0);
    io_sharedInputs_0_arw_payload_len : in unsigned(7 downto 0);
    io_sharedInputs_0_arw_payload_size : in unsigned(2 downto 0);
    io_sharedInputs_0_arw_payload_burst : in std_logic_vector(1 downto 0);
    io_sharedInputs_0_arw_payload_write : in std_logic;
    io_sharedInputs_0_w_valid : in std_logic;
    io_sharedInputs_0_w_ready : out std_logic;
    io_sharedInputs_0_w_payload_data : in std_logic_vector(31 downto 0);
    io_sharedInputs_0_w_payload_strb : in std_logic_vector(3 downto 0);
    io_sharedInputs_0_w_payload_last : in std_logic;
    io_sharedInputs_0_b_valid : out std_logic;
    io_sharedInputs_0_b_ready : in std_logic;
    io_sharedInputs_0_b_payload_id : out unsigned(2 downto 0);
    io_sharedInputs_0_b_payload_resp : out std_logic_vector(1 downto 0);
    io_sharedInputs_0_r_valid : out std_logic;
    io_sharedInputs_0_r_ready : in std_logic;
    io_sharedInputs_0_r_payload_data : out std_logic_vector(31 downto 0);
    io_sharedInputs_0_r_payload_id : out unsigned(2 downto 0);
    io_sharedInputs_0_r_payload_resp : out std_logic_vector(1 downto 0);
    io_sharedInputs_0_r_payload_last : out std_logic;
    io_output_arw_valid : out std_logic;
    io_output_arw_ready : in std_logic;
    io_output_arw_payload_addr : out unsigned(14 downto 0);
    io_output_arw_payload_id : out unsigned(3 downto 0);
    io_output_arw_payload_len : out unsigned(7 downto 0);
    io_output_arw_payload_size : out unsigned(2 downto 0);
    io_output_arw_payload_burst : out std_logic_vector(1 downto 0);
    io_output_arw_payload_write : out std_logic;
    io_output_w_valid : out std_logic;
    io_output_w_ready : in std_logic;
    io_output_w_payload_data : out std_logic_vector(31 downto 0);
    io_output_w_payload_strb : out std_logic_vector(3 downto 0);
    io_output_w_payload_last : out std_logic;
    io_output_b_valid : in std_logic;
    io_output_b_ready : out std_logic;
    io_output_b_payload_id : in unsigned(3 downto 0);
    io_output_b_payload_resp : in std_logic_vector(1 downto 0);
    io_output_r_valid : in std_logic;
    io_output_r_ready : out std_logic;
    io_output_r_payload_data : in std_logic_vector(31 downto 0);
    io_output_r_payload_id : in unsigned(3 downto 0);
    io_output_r_payload_resp : in std_logic_vector(1 downto 0);
    io_output_r_payload_last : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4SharedArbiter;

architecture arch of Axi4SharedArbiter is
  signal cmdArbiter_io_output_fork_io_outputs_1_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_ready : std_logic;
  signal io_sharedInputs_0_w_ready_read_buffer : std_logic;
  signal io_output_w_valid_read_buffer : std_logic;
  signal io_output_w_payload_last_read_buffer : std_logic;
  signal cmdArbiter_io_inputs_0_ready : std_logic;
  signal cmdArbiter_io_inputs_1_ready : std_logic;
  signal cmdArbiter_io_output_valid : std_logic;
  signal cmdArbiter_io_output_payload_addr : unsigned(14 downto 0);
  signal cmdArbiter_io_output_payload_id : unsigned(2 downto 0);
  signal cmdArbiter_io_output_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_payload_write : std_logic;
  signal cmdArbiter_io_chosen : unsigned(0 downto 0);
  signal cmdArbiter_io_chosenOH : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_input_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_0_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_addr : unsigned(14 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_id : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_write : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_addr : unsigned(14 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_id : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_write : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_push_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_occupancy : unsigned(2 downto 0);
  signal zz_io_output_r_ready : std_logic;

  signal inputsCmd_0_valid : std_logic;
  signal inputsCmd_0_ready : std_logic;
  signal inputsCmd_0_payload_addr : unsigned(14 downto 0);
  signal inputsCmd_0_payload_id : unsigned(2 downto 0);
  signal inputsCmd_0_payload_len : unsigned(7 downto 0);
  signal inputsCmd_0_payload_size : unsigned(2 downto 0);
  signal inputsCmd_0_payload_burst : std_logic_vector(1 downto 0);
  signal inputsCmd_0_payload_write : std_logic;
  signal inputsCmd_1_valid : std_logic;
  signal inputsCmd_1_ready : std_logic;
  signal inputsCmd_1_payload_addr : unsigned(14 downto 0);
  signal inputsCmd_1_payload_id : unsigned(2 downto 0);
  signal inputsCmd_1_payload_len : unsigned(7 downto 0);
  signal inputsCmd_1_payload_size : unsigned(2 downto 0);
  signal inputsCmd_1_payload_burst : std_logic_vector(1 downto 0);
  signal inputsCmd_1_payload_write : std_logic;
  signal zz_io_output_arw_payload_id : std_logic;
  signal when_Stream_l408 : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_addr : unsigned(14 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_id : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_write : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_ready : std_logic;
  signal writeLogic_routeDataInput_valid : std_logic;
  signal writeLogic_routeDataInput_ready : std_logic;
  signal writeLogic_routeDataInput_payload_data : std_logic_vector(31 downto 0);
  signal writeLogic_routeDataInput_payload_strb : std_logic_vector(3 downto 0);
  signal writeLogic_routeDataInput_payload_last : std_logic;
  signal io_output_w_fire : std_logic;
  signal writeLogic_writeRspSels_0 : std_logic;
  signal readRspIndex : unsigned(0 downto 0);
  signal readRspSels_0 : std_logic;
  signal readRspSels_1 : std_logic;
begin
  io_sharedInputs_0_w_ready <= io_sharedInputs_0_w_ready_read_buffer;
  io_output_w_valid <= io_output_w_valid_read_buffer;
  io_output_w_payload_last <= io_output_w_payload_last_read_buffer;
  cmdArbiter : entity work.StreamArbiter
    port map ( 
      io_inputs_0_valid => inputsCmd_0_valid,
      io_inputs_0_ready => cmdArbiter_io_inputs_0_ready,
      io_inputs_0_payload_addr => inputsCmd_0_payload_addr,
      io_inputs_0_payload_id => inputsCmd_0_payload_id,
      io_inputs_0_payload_len => inputsCmd_0_payload_len,
      io_inputs_0_payload_size => inputsCmd_0_payload_size,
      io_inputs_0_payload_burst => inputsCmd_0_payload_burst,
      io_inputs_0_payload_write => inputsCmd_0_payload_write,
      io_inputs_1_valid => inputsCmd_1_valid,
      io_inputs_1_ready => cmdArbiter_io_inputs_1_ready,
      io_inputs_1_payload_addr => inputsCmd_1_payload_addr,
      io_inputs_1_payload_id => inputsCmd_1_payload_id,
      io_inputs_1_payload_len => inputsCmd_1_payload_len,
      io_inputs_1_payload_size => inputsCmd_1_payload_size,
      io_inputs_1_payload_burst => inputsCmd_1_payload_burst,
      io_inputs_1_payload_write => inputsCmd_1_payload_write,
      io_output_valid => cmdArbiter_io_output_valid,
      io_output_ready => cmdArbiter_io_output_fork_io_input_ready,
      io_output_payload_addr => cmdArbiter_io_output_payload_addr,
      io_output_payload_id => cmdArbiter_io_output_payload_id,
      io_output_payload_len => cmdArbiter_io_output_payload_len,
      io_output_payload_size => cmdArbiter_io_output_payload_size,
      io_output_payload_burst => cmdArbiter_io_output_payload_burst,
      io_output_payload_write => cmdArbiter_io_output_payload_write,
      io_chosen => cmdArbiter_io_chosen,
      io_chosenOH => cmdArbiter_io_chosenOH,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  cmdArbiter_io_output_fork : entity work.StreamFork
    port map ( 
      io_input_valid => cmdArbiter_io_output_valid,
      io_input_ready => cmdArbiter_io_output_fork_io_input_ready,
      io_input_payload_addr => cmdArbiter_io_output_payload_addr,
      io_input_payload_id => cmdArbiter_io_output_payload_id,
      io_input_payload_len => cmdArbiter_io_output_payload_len,
      io_input_payload_size => cmdArbiter_io_output_payload_size,
      io_input_payload_burst => cmdArbiter_io_output_payload_burst,
      io_input_payload_write => cmdArbiter_io_output_payload_write,
      io_outputs_0_valid => cmdArbiter_io_output_fork_io_outputs_0_valid,
      io_outputs_0_ready => io_output_arw_ready,
      io_outputs_0_payload_addr => cmdArbiter_io_output_fork_io_outputs_0_payload_addr,
      io_outputs_0_payload_id => cmdArbiter_io_output_fork_io_outputs_0_payload_id,
      io_outputs_0_payload_len => cmdArbiter_io_output_fork_io_outputs_0_payload_len,
      io_outputs_0_payload_size => cmdArbiter_io_output_fork_io_outputs_0_payload_size,
      io_outputs_0_payload_burst => cmdArbiter_io_output_fork_io_outputs_0_payload_burst,
      io_outputs_0_payload_write => cmdArbiter_io_output_fork_io_outputs_0_payload_write,
      io_outputs_1_valid => cmdArbiter_io_output_fork_io_outputs_1_valid,
      io_outputs_1_ready => cmdArbiter_io_output_fork_io_outputs_1_ready,
      io_outputs_1_payload_addr => cmdArbiter_io_output_fork_io_outputs_1_payload_addr,
      io_outputs_1_payload_id => cmdArbiter_io_output_fork_io_outputs_1_payload_id,
      io_outputs_1_payload_len => cmdArbiter_io_output_fork_io_outputs_1_payload_len,
      io_outputs_1_payload_size => cmdArbiter_io_output_fork_io_outputs_1_payload_size,
      io_outputs_1_payload_burst => cmdArbiter_io_output_fork_io_outputs_1_payload_burst,
      io_outputs_1_payload_write => cmdArbiter_io_output_fork_io_outputs_1_payload_write,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo : entity work.StreamFifoLowLatency
    port map ( 
      io_push_valid => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_valid,
      io_push_ready => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_push_ready,
      io_pop_valid => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid,
      io_pop_ready => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_ready,
      io_flush => pkg_toStdLogic(false),
      io_occupancy => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_occupancy,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  process(readRspIndex,io_readInputs_0_r_ready,io_sharedInputs_0_r_ready)
  begin
    case readRspIndex is
      when "0" =>
        zz_io_output_r_ready <= io_readInputs_0_r_ready;
      when others =>
        zz_io_output_r_ready <= io_sharedInputs_0_r_ready;
    end case;
  end process;

  inputsCmd_0_valid <= io_readInputs_0_ar_valid;
  io_readInputs_0_ar_ready <= inputsCmd_0_ready;
  inputsCmd_0_payload_addr <= io_readInputs_0_ar_payload_addr;
  inputsCmd_0_payload_id <= io_readInputs_0_ar_payload_id;
  inputsCmd_0_payload_len <= io_readInputs_0_ar_payload_len;
  inputsCmd_0_payload_size <= io_readInputs_0_ar_payload_size;
  inputsCmd_0_payload_burst <= io_readInputs_0_ar_payload_burst;
  inputsCmd_0_payload_write <= pkg_toStdLogic(false);
  inputsCmd_1_valid <= io_sharedInputs_0_arw_valid;
  io_sharedInputs_0_arw_ready <= inputsCmd_1_ready;
  inputsCmd_1_payload_addr <= io_sharedInputs_0_arw_payload_addr;
  inputsCmd_1_payload_id <= io_sharedInputs_0_arw_payload_id;
  inputsCmd_1_payload_len <= io_sharedInputs_0_arw_payload_len;
  inputsCmd_1_payload_size <= io_sharedInputs_0_arw_payload_size;
  inputsCmd_1_payload_burst <= io_sharedInputs_0_arw_payload_burst;
  inputsCmd_1_payload_write <= io_sharedInputs_0_arw_payload_write;
  inputsCmd_0_ready <= cmdArbiter_io_inputs_0_ready;
  inputsCmd_1_ready <= cmdArbiter_io_inputs_1_ready;
  io_output_arw_valid <= cmdArbiter_io_output_fork_io_outputs_0_valid;
  io_output_arw_payload_addr <= cmdArbiter_io_output_fork_io_outputs_0_payload_addr;
  io_output_arw_payload_len <= cmdArbiter_io_output_fork_io_outputs_0_payload_len;
  io_output_arw_payload_size <= cmdArbiter_io_output_fork_io_outputs_0_payload_size;
  io_output_arw_payload_burst <= cmdArbiter_io_output_fork_io_outputs_0_payload_burst;
  io_output_arw_payload_write <= cmdArbiter_io_output_fork_io_outputs_0_payload_write;
  zz_io_output_arw_payload_id <= pkg_extract(pkg_cat(pkg_extract(cmdArbiter_io_chosenOH,1,1),pkg_extract(cmdArbiter_io_chosenOH,0,0)),1);
  io_output_arw_payload_id <= pkg_mux(cmdArbiter_io_output_fork_io_outputs_0_payload_write,pkg_resize(unsigned(std_logic_vector(cmdArbiter_io_output_fork_io_outputs_0_payload_id)),4),unsigned(pkg_cat(std_logic_vector(unsigned(pkg_toStdLogicVector(zz_io_output_arw_payload_id))),std_logic_vector(cmdArbiter_io_output_fork_io_outputs_0_payload_id))));
  when_Stream_l408 <= (not cmdArbiter_io_output_fork_io_outputs_1_payload_write);
  process(cmdArbiter_io_output_fork_io_outputs_1_valid,when_Stream_l408)
  begin
    cmdArbiter_io_output_fork_io_outputs_1_thrown_valid <= cmdArbiter_io_output_fork_io_outputs_1_valid;
    if when_Stream_l408 = '1' then
      cmdArbiter_io_output_fork_io_outputs_1_thrown_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  process(cmdArbiter_io_output_fork_io_outputs_1_thrown_ready,when_Stream_l408)
  begin
    cmdArbiter_io_output_fork_io_outputs_1_ready <= cmdArbiter_io_output_fork_io_outputs_1_thrown_ready;
    if when_Stream_l408 = '1' then
      cmdArbiter_io_output_fork_io_outputs_1_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_addr <= cmdArbiter_io_output_fork_io_outputs_1_payload_addr;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_id <= cmdArbiter_io_output_fork_io_outputs_1_payload_id;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_len <= cmdArbiter_io_output_fork_io_outputs_1_payload_len;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_size <= cmdArbiter_io_output_fork_io_outputs_1_payload_size;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_burst <= cmdArbiter_io_output_fork_io_outputs_1_payload_burst;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_write <= cmdArbiter_io_output_fork_io_outputs_1_payload_write;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_valid <= cmdArbiter_io_output_fork_io_outputs_1_thrown_valid;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_ready <= cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_ready;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_ready <= cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_push_ready;
  writeLogic_routeDataInput_valid <= io_sharedInputs_0_w_valid;
  writeLogic_routeDataInput_ready <= io_sharedInputs_0_w_ready_read_buffer;
  writeLogic_routeDataInput_payload_data <= io_sharedInputs_0_w_payload_data;
  writeLogic_routeDataInput_payload_strb <= io_sharedInputs_0_w_payload_strb;
  writeLogic_routeDataInput_payload_last <= io_sharedInputs_0_w_payload_last;
  io_output_w_valid_read_buffer <= (cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid and writeLogic_routeDataInput_valid);
  io_output_w_payload_data <= writeLogic_routeDataInput_payload_data;
  io_output_w_payload_strb <= writeLogic_routeDataInput_payload_strb;
  io_output_w_payload_last_read_buffer <= writeLogic_routeDataInput_payload_last;
  io_sharedInputs_0_w_ready_read_buffer <= ((cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid and io_output_w_ready) and pkg_toStdLogic(true));
  io_output_w_fire <= (io_output_w_valid_read_buffer and io_output_w_ready);
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_ready <= (io_output_w_fire and io_output_w_payload_last_read_buffer);
  writeLogic_writeRspSels_0 <= pkg_toStdLogic(true);
  io_sharedInputs_0_b_valid <= (io_output_b_valid and writeLogic_writeRspSels_0);
  io_sharedInputs_0_b_payload_resp <= io_output_b_payload_resp;
  io_sharedInputs_0_b_payload_id <= pkg_resize(io_output_b_payload_id,3);
  io_output_b_ready <= io_sharedInputs_0_b_ready;
  readRspIndex <= pkg_extract(io_output_r_payload_id,3,3);
  readRspSels_0 <= pkg_toStdLogic(readRspIndex = pkg_unsigned("0"));
  readRspSels_1 <= pkg_toStdLogic(readRspIndex = pkg_unsigned("1"));
  io_readInputs_0_r_valid <= (io_output_r_valid and readRspSels_0);
  io_readInputs_0_r_payload_data <= io_output_r_payload_data;
  io_readInputs_0_r_payload_resp <= io_output_r_payload_resp;
  io_readInputs_0_r_payload_last <= io_output_r_payload_last;
  io_readInputs_0_r_payload_id <= pkg_resize(io_output_r_payload_id,3);
  io_sharedInputs_0_r_valid <= (io_output_r_valid and readRspSels_1);
  io_sharedInputs_0_r_payload_data <= io_output_r_payload_data;
  io_sharedInputs_0_r_payload_resp <= io_output_r_payload_resp;
  io_sharedInputs_0_r_payload_last <= io_output_r_payload_last;
  io_sharedInputs_0_r_payload_id <= pkg_resize(io_output_r_payload_id,3);
  io_output_r_ready <= zz_io_output_r_ready;
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Axi4SharedArbiter_1 is
  port(
    io_sharedInputs_0_arw_valid : in std_logic;
    io_sharedInputs_0_arw_ready : out std_logic;
    io_sharedInputs_0_arw_payload_addr : in unsigned(19 downto 0);
    io_sharedInputs_0_arw_payload_id : in unsigned(3 downto 0);
    io_sharedInputs_0_arw_payload_len : in unsigned(7 downto 0);
    io_sharedInputs_0_arw_payload_size : in unsigned(2 downto 0);
    io_sharedInputs_0_arw_payload_burst : in std_logic_vector(1 downto 0);
    io_sharedInputs_0_arw_payload_write : in std_logic;
    io_sharedInputs_0_w_valid : in std_logic;
    io_sharedInputs_0_w_ready : out std_logic;
    io_sharedInputs_0_w_payload_data : in std_logic_vector(31 downto 0);
    io_sharedInputs_0_w_payload_strb : in std_logic_vector(3 downto 0);
    io_sharedInputs_0_w_payload_last : in std_logic;
    io_sharedInputs_0_b_valid : out std_logic;
    io_sharedInputs_0_b_ready : in std_logic;
    io_sharedInputs_0_b_payload_id : out unsigned(3 downto 0);
    io_sharedInputs_0_b_payload_resp : out std_logic_vector(1 downto 0);
    io_sharedInputs_0_r_valid : out std_logic;
    io_sharedInputs_0_r_ready : in std_logic;
    io_sharedInputs_0_r_payload_data : out std_logic_vector(31 downto 0);
    io_sharedInputs_0_r_payload_id : out unsigned(3 downto 0);
    io_sharedInputs_0_r_payload_resp : out std_logic_vector(1 downto 0);
    io_sharedInputs_0_r_payload_last : out std_logic;
    io_output_arw_valid : out std_logic;
    io_output_arw_ready : in std_logic;
    io_output_arw_payload_addr : out unsigned(19 downto 0);
    io_output_arw_payload_id : out unsigned(3 downto 0);
    io_output_arw_payload_len : out unsigned(7 downto 0);
    io_output_arw_payload_size : out unsigned(2 downto 0);
    io_output_arw_payload_burst : out std_logic_vector(1 downto 0);
    io_output_arw_payload_write : out std_logic;
    io_output_w_valid : out std_logic;
    io_output_w_ready : in std_logic;
    io_output_w_payload_data : out std_logic_vector(31 downto 0);
    io_output_w_payload_strb : out std_logic_vector(3 downto 0);
    io_output_w_payload_last : out std_logic;
    io_output_b_valid : in std_logic;
    io_output_b_ready : out std_logic;
    io_output_b_payload_id : in unsigned(3 downto 0);
    io_output_b_payload_resp : in std_logic_vector(1 downto 0);
    io_output_r_valid : in std_logic;
    io_output_r_ready : out std_logic;
    io_output_r_payload_data : in std_logic_vector(31 downto 0);
    io_output_r_payload_id : in unsigned(3 downto 0);
    io_output_r_payload_resp : in std_logic_vector(1 downto 0);
    io_output_r_payload_last : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Axi4SharedArbiter_1;

architecture arch of Axi4SharedArbiter_1 is
  signal cmdArbiter_io_output_fork_io_outputs_1_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_ready : std_logic;
  signal io_sharedInputs_0_w_ready_read_buffer : std_logic;
  signal io_output_w_valid_read_buffer : std_logic;
  signal io_output_w_payload_last_read_buffer : std_logic;
  signal cmdArbiter_io_inputs_0_ready : std_logic;
  signal cmdArbiter_io_output_valid : std_logic;
  signal cmdArbiter_io_output_payload_addr : unsigned(19 downto 0);
  signal cmdArbiter_io_output_payload_id : unsigned(3 downto 0);
  signal cmdArbiter_io_output_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_payload_write : std_logic;
  signal cmdArbiter_io_chosenOH : std_logic_vector(0 downto 0);
  signal cmdArbiter_io_output_fork_io_input_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_0_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_addr : unsigned(19 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_id : unsigned(3 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_0_payload_write : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_addr : unsigned(19 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_id : unsigned(3 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_payload_write : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_push_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_occupancy : unsigned(2 downto 0);

  signal inputsCmd_0_valid : std_logic;
  signal inputsCmd_0_ready : std_logic;
  signal inputsCmd_0_payload_addr : unsigned(19 downto 0);
  signal inputsCmd_0_payload_id : unsigned(3 downto 0);
  signal inputsCmd_0_payload_len : unsigned(7 downto 0);
  signal inputsCmd_0_payload_size : unsigned(2 downto 0);
  signal inputsCmd_0_payload_burst : std_logic_vector(1 downto 0);
  signal inputsCmd_0_payload_write : std_logic;
  signal when_Stream_l408 : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_ready : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_addr : unsigned(19 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_id : unsigned(3 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_len : unsigned(7 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_size : unsigned(2 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_burst : std_logic_vector(1 downto 0);
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_write : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_valid : std_logic;
  signal cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_ready : std_logic;
  signal writeLogic_routeDataInput_valid : std_logic;
  signal writeLogic_routeDataInput_ready : std_logic;
  signal writeLogic_routeDataInput_payload_data : std_logic_vector(31 downto 0);
  signal writeLogic_routeDataInput_payload_strb : std_logic_vector(3 downto 0);
  signal writeLogic_routeDataInput_payload_last : std_logic;
  signal io_output_w_fire : std_logic;
  signal writeLogic_writeRspSels_0 : std_logic;
  signal readRspSels_0 : std_logic;
begin
  io_sharedInputs_0_w_ready <= io_sharedInputs_0_w_ready_read_buffer;
  io_output_w_valid <= io_output_w_valid_read_buffer;
  io_output_w_payload_last <= io_output_w_payload_last_read_buffer;
  cmdArbiter : entity work.StreamArbiter_1
    port map ( 
      io_inputs_0_valid => inputsCmd_0_valid,
      io_inputs_0_ready => cmdArbiter_io_inputs_0_ready,
      io_inputs_0_payload_addr => inputsCmd_0_payload_addr,
      io_inputs_0_payload_id => inputsCmd_0_payload_id,
      io_inputs_0_payload_len => inputsCmd_0_payload_len,
      io_inputs_0_payload_size => inputsCmd_0_payload_size,
      io_inputs_0_payload_burst => inputsCmd_0_payload_burst,
      io_inputs_0_payload_write => inputsCmd_0_payload_write,
      io_output_valid => cmdArbiter_io_output_valid,
      io_output_ready => cmdArbiter_io_output_fork_io_input_ready,
      io_output_payload_addr => cmdArbiter_io_output_payload_addr,
      io_output_payload_id => cmdArbiter_io_output_payload_id,
      io_output_payload_len => cmdArbiter_io_output_payload_len,
      io_output_payload_size => cmdArbiter_io_output_payload_size,
      io_output_payload_burst => cmdArbiter_io_output_payload_burst,
      io_output_payload_write => cmdArbiter_io_output_payload_write,
      io_chosenOH => cmdArbiter_io_chosenOH,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  cmdArbiter_io_output_fork : entity work.StreamFork_1
    port map ( 
      io_input_valid => cmdArbiter_io_output_valid,
      io_input_ready => cmdArbiter_io_output_fork_io_input_ready,
      io_input_payload_addr => cmdArbiter_io_output_payload_addr,
      io_input_payload_id => cmdArbiter_io_output_payload_id,
      io_input_payload_len => cmdArbiter_io_output_payload_len,
      io_input_payload_size => cmdArbiter_io_output_payload_size,
      io_input_payload_burst => cmdArbiter_io_output_payload_burst,
      io_input_payload_write => cmdArbiter_io_output_payload_write,
      io_outputs_0_valid => cmdArbiter_io_output_fork_io_outputs_0_valid,
      io_outputs_0_ready => io_output_arw_ready,
      io_outputs_0_payload_addr => cmdArbiter_io_output_fork_io_outputs_0_payload_addr,
      io_outputs_0_payload_id => cmdArbiter_io_output_fork_io_outputs_0_payload_id,
      io_outputs_0_payload_len => cmdArbiter_io_output_fork_io_outputs_0_payload_len,
      io_outputs_0_payload_size => cmdArbiter_io_output_fork_io_outputs_0_payload_size,
      io_outputs_0_payload_burst => cmdArbiter_io_output_fork_io_outputs_0_payload_burst,
      io_outputs_0_payload_write => cmdArbiter_io_output_fork_io_outputs_0_payload_write,
      io_outputs_1_valid => cmdArbiter_io_output_fork_io_outputs_1_valid,
      io_outputs_1_ready => cmdArbiter_io_output_fork_io_outputs_1_ready,
      io_outputs_1_payload_addr => cmdArbiter_io_output_fork_io_outputs_1_payload_addr,
      io_outputs_1_payload_id => cmdArbiter_io_output_fork_io_outputs_1_payload_id,
      io_outputs_1_payload_len => cmdArbiter_io_output_fork_io_outputs_1_payload_len,
      io_outputs_1_payload_size => cmdArbiter_io_output_fork_io_outputs_1_payload_size,
      io_outputs_1_payload_burst => cmdArbiter_io_output_fork_io_outputs_1_payload_burst,
      io_outputs_1_payload_write => cmdArbiter_io_output_fork_io_outputs_1_payload_write,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo : entity work.StreamFifoLowLatency
    port map ( 
      io_push_valid => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_valid,
      io_push_ready => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_push_ready,
      io_pop_valid => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid,
      io_pop_ready => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_ready,
      io_flush => pkg_toStdLogic(false),
      io_occupancy => cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_occupancy,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  inputsCmd_0_valid <= io_sharedInputs_0_arw_valid;
  io_sharedInputs_0_arw_ready <= inputsCmd_0_ready;
  inputsCmd_0_payload_addr <= io_sharedInputs_0_arw_payload_addr;
  inputsCmd_0_payload_id <= io_sharedInputs_0_arw_payload_id;
  inputsCmd_0_payload_len <= io_sharedInputs_0_arw_payload_len;
  inputsCmd_0_payload_size <= io_sharedInputs_0_arw_payload_size;
  inputsCmd_0_payload_burst <= io_sharedInputs_0_arw_payload_burst;
  inputsCmd_0_payload_write <= io_sharedInputs_0_arw_payload_write;
  inputsCmd_0_ready <= cmdArbiter_io_inputs_0_ready;
  io_output_arw_valid <= cmdArbiter_io_output_fork_io_outputs_0_valid;
  io_output_arw_payload_addr <= cmdArbiter_io_output_fork_io_outputs_0_payload_addr;
  io_output_arw_payload_len <= cmdArbiter_io_output_fork_io_outputs_0_payload_len;
  io_output_arw_payload_size <= cmdArbiter_io_output_fork_io_outputs_0_payload_size;
  io_output_arw_payload_burst <= cmdArbiter_io_output_fork_io_outputs_0_payload_burst;
  io_output_arw_payload_write <= cmdArbiter_io_output_fork_io_outputs_0_payload_write;
  io_output_arw_payload_id <= pkg_mux(cmdArbiter_io_output_fork_io_outputs_0_payload_write,unsigned(std_logic_vector(cmdArbiter_io_output_fork_io_outputs_0_payload_id)),unsigned(std_logic_vector(cmdArbiter_io_output_fork_io_outputs_0_payload_id)));
  when_Stream_l408 <= (not cmdArbiter_io_output_fork_io_outputs_1_payload_write);
  process(cmdArbiter_io_output_fork_io_outputs_1_valid,when_Stream_l408)
  begin
    cmdArbiter_io_output_fork_io_outputs_1_thrown_valid <= cmdArbiter_io_output_fork_io_outputs_1_valid;
    if when_Stream_l408 = '1' then
      cmdArbiter_io_output_fork_io_outputs_1_thrown_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  process(cmdArbiter_io_output_fork_io_outputs_1_thrown_ready,when_Stream_l408)
  begin
    cmdArbiter_io_output_fork_io_outputs_1_ready <= cmdArbiter_io_output_fork_io_outputs_1_thrown_ready;
    if when_Stream_l408 = '1' then
      cmdArbiter_io_output_fork_io_outputs_1_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_addr <= cmdArbiter_io_output_fork_io_outputs_1_payload_addr;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_id <= cmdArbiter_io_output_fork_io_outputs_1_payload_id;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_len <= cmdArbiter_io_output_fork_io_outputs_1_payload_len;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_size <= cmdArbiter_io_output_fork_io_outputs_1_payload_size;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_burst <= cmdArbiter_io_output_fork_io_outputs_1_payload_burst;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_payload_write <= cmdArbiter_io_output_fork_io_outputs_1_payload_write;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_valid <= cmdArbiter_io_output_fork_io_outputs_1_thrown_valid;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_ready <= cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_ready;
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_ready <= cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_push_ready;
  writeLogic_routeDataInput_valid <= io_sharedInputs_0_w_valid;
  writeLogic_routeDataInput_ready <= io_sharedInputs_0_w_ready_read_buffer;
  writeLogic_routeDataInput_payload_data <= io_sharedInputs_0_w_payload_data;
  writeLogic_routeDataInput_payload_strb <= io_sharedInputs_0_w_payload_strb;
  writeLogic_routeDataInput_payload_last <= io_sharedInputs_0_w_payload_last;
  io_output_w_valid_read_buffer <= (cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid and writeLogic_routeDataInput_valid);
  io_output_w_payload_data <= writeLogic_routeDataInput_payload_data;
  io_output_w_payload_strb <= writeLogic_routeDataInput_payload_strb;
  io_output_w_payload_last_read_buffer <= writeLogic_routeDataInput_payload_last;
  io_sharedInputs_0_w_ready_read_buffer <= ((cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_valid and io_output_w_ready) and pkg_toStdLogic(true));
  io_output_w_fire <= (io_output_w_valid_read_buffer and io_output_w_ready);
  cmdArbiter_io_output_fork_io_outputs_1_thrown_translated_fifo_io_pop_ready <= (io_output_w_fire and io_output_w_payload_last_read_buffer);
  writeLogic_writeRspSels_0 <= pkg_toStdLogic(true);
  io_sharedInputs_0_b_valid <= (io_output_b_valid and writeLogic_writeRspSels_0);
  io_sharedInputs_0_b_payload_resp <= io_output_b_payload_resp;
  io_sharedInputs_0_b_payload_id <= io_output_b_payload_id;
  io_output_b_ready <= io_sharedInputs_0_b_ready;
  readRspSels_0 <= pkg_toStdLogic(true);
  io_sharedInputs_0_r_valid <= (io_output_r_valid and readRspSels_0);
  io_sharedInputs_0_r_payload_data <= io_output_r_payload_data;
  io_sharedInputs_0_r_payload_resp <= io_output_r_payload_resp;
  io_sharedInputs_0_r_payload_last <= io_output_r_payload_last;
  io_sharedInputs_0_r_payload_id <= io_output_r_payload_id;
  io_output_r_ready <= io_sharedInputs_0_r_ready;
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Apb3Decoder is
  port(
    io_input_PADDR : in unsigned(19 downto 0);
    io_input_PSEL : in std_logic_vector(0 downto 0);
    io_input_PENABLE : in std_logic;
    io_input_PREADY : out std_logic;
    io_input_PWRITE : in std_logic;
    io_input_PWDATA : in std_logic_vector(31 downto 0);
    io_input_PRDATA : out std_logic_vector(31 downto 0);
    io_input_PSLVERROR : out std_logic;
    io_output_PADDR : out unsigned(19 downto 0);
    io_output_PSEL : out std_logic_vector(2 downto 0);
    io_output_PENABLE : out std_logic;
    io_output_PREADY : in std_logic;
    io_output_PWRITE : out std_logic;
    io_output_PWDATA : out std_logic_vector(31 downto 0);
    io_output_PRDATA : in std_logic_vector(31 downto 0);
    io_output_PSLVERROR : in std_logic
  );
end Apb3Decoder;

architecture arch of Apb3Decoder is
  signal io_output_PSEL_read_buffer : std_logic_vector(2 downto 0);

  signal when_Apb3Decoder_l88 : std_logic;
begin
  io_output_PSEL <= io_output_PSEL_read_buffer;
  io_output_PADDR <= io_input_PADDR;
  io_output_PENABLE <= io_input_PENABLE;
  io_output_PWRITE <= io_input_PWRITE;
  io_output_PWDATA <= io_input_PWDATA;
  process(io_input_PADDR,io_input_PSEL)
  begin
    io_output_PSEL_read_buffer(0) <= (pkg_toStdLogic((io_input_PADDR and pkg_not(pkg_unsigned("00000000111111111111"))) = pkg_unsigned("00000000000000000000")) and pkg_extract(io_input_PSEL,0));
    io_output_PSEL_read_buffer(1) <= (pkg_toStdLogic((io_input_PADDR and pkg_not(pkg_unsigned("00000000111111111111"))) = pkg_unsigned("00010000000000000000")) and pkg_extract(io_input_PSEL,0));
    io_output_PSEL_read_buffer(2) <= (pkg_toStdLogic((io_input_PADDR and pkg_not(pkg_unsigned("00000000111111111111"))) = pkg_unsigned("00100000000000000000")) and pkg_extract(io_input_PSEL,0));
  end process;

  process(io_output_PREADY,when_Apb3Decoder_l88)
  begin
    io_input_PREADY <= io_output_PREADY;
    if when_Apb3Decoder_l88 = '1' then
      io_input_PREADY <= pkg_toStdLogic(true);
    end if;
  end process;

  io_input_PRDATA <= io_output_PRDATA;
  process(io_output_PSLVERROR,when_Apb3Decoder_l88)
  begin
    io_input_PSLVERROR <= io_output_PSLVERROR;
    if when_Apb3Decoder_l88 = '1' then
      io_input_PSLVERROR <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Apb3Decoder_l88 <= (pkg_extract(io_input_PSEL,0) and pkg_toStdLogic(io_output_PSEL_read_buffer = pkg_stdLogicVector("000")));
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Apb3Router is
  port(
    io_input_PADDR : in unsigned(19 downto 0);
    io_input_PSEL : in std_logic_vector(2 downto 0);
    io_input_PENABLE : in std_logic;
    io_input_PREADY : out std_logic;
    io_input_PWRITE : in std_logic;
    io_input_PWDATA : in std_logic_vector(31 downto 0);
    io_input_PRDATA : out std_logic_vector(31 downto 0);
    io_input_PSLVERROR : out std_logic;
    io_outputs_0_PADDR : out unsigned(19 downto 0);
    io_outputs_0_PSEL : out std_logic_vector(0 downto 0);
    io_outputs_0_PENABLE : out std_logic;
    io_outputs_0_PREADY : in std_logic;
    io_outputs_0_PWRITE : out std_logic;
    io_outputs_0_PWDATA : out std_logic_vector(31 downto 0);
    io_outputs_0_PRDATA : in std_logic_vector(31 downto 0);
    io_outputs_0_PSLVERROR : in std_logic;
    io_outputs_1_PADDR : out unsigned(19 downto 0);
    io_outputs_1_PSEL : out std_logic_vector(0 downto 0);
    io_outputs_1_PENABLE : out std_logic;
    io_outputs_1_PREADY : in std_logic;
    io_outputs_1_PWRITE : out std_logic;
    io_outputs_1_PWDATA : out std_logic_vector(31 downto 0);
    io_outputs_1_PRDATA : in std_logic_vector(31 downto 0);
    io_outputs_1_PSLVERROR : in std_logic;
    io_outputs_2_PADDR : out unsigned(19 downto 0);
    io_outputs_2_PSEL : out std_logic_vector(0 downto 0);
    io_outputs_2_PENABLE : out std_logic;
    io_outputs_2_PREADY : in std_logic;
    io_outputs_2_PWRITE : out std_logic;
    io_outputs_2_PWDATA : out std_logic_vector(31 downto 0);
    io_outputs_2_PRDATA : in std_logic_vector(31 downto 0);
    io_outputs_2_PSLVERROR : in std_logic;
    io_mainClk : in std_logic;
    resetCtrl_axiReset : in std_logic
  );
end Apb3Router;

architecture arch of Apb3Router is
  signal zz_io_input_PREADY : std_logic;
  signal zz_io_input_PRDATA : std_logic_vector(31 downto 0);
  signal zz_io_input_PSLVERROR : std_logic;

  signal zz_selIndex : std_logic;
  signal zz_selIndex_1 : std_logic;
  signal selIndex : unsigned(1 downto 0);
begin
  process(selIndex,io_outputs_0_PREADY,io_outputs_0_PRDATA,io_outputs_0_PSLVERROR,io_outputs_1_PREADY,io_outputs_1_PRDATA,io_outputs_1_PSLVERROR,io_outputs_2_PREADY,io_outputs_2_PRDATA,io_outputs_2_PSLVERROR)
  begin
    case selIndex is
      when "00" =>
        zz_io_input_PREADY <= io_outputs_0_PREADY;
        zz_io_input_PRDATA <= io_outputs_0_PRDATA;
        zz_io_input_PSLVERROR <= io_outputs_0_PSLVERROR;
      when "01" =>
        zz_io_input_PREADY <= io_outputs_1_PREADY;
        zz_io_input_PRDATA <= io_outputs_1_PRDATA;
        zz_io_input_PSLVERROR <= io_outputs_1_PSLVERROR;
      when others =>
        zz_io_input_PREADY <= io_outputs_2_PREADY;
        zz_io_input_PRDATA <= io_outputs_2_PRDATA;
        zz_io_input_PSLVERROR <= io_outputs_2_PSLVERROR;
    end case;
  end process;

  io_outputs_0_PADDR <= io_input_PADDR;
  io_outputs_0_PENABLE <= io_input_PENABLE;
  io_outputs_0_PSEL(0) <= pkg_extract(io_input_PSEL,0);
  io_outputs_0_PWRITE <= io_input_PWRITE;
  io_outputs_0_PWDATA <= io_input_PWDATA;
  io_outputs_1_PADDR <= io_input_PADDR;
  io_outputs_1_PENABLE <= io_input_PENABLE;
  io_outputs_1_PSEL(0) <= pkg_extract(io_input_PSEL,1);
  io_outputs_1_PWRITE <= io_input_PWRITE;
  io_outputs_1_PWDATA <= io_input_PWDATA;
  io_outputs_2_PADDR <= io_input_PADDR;
  io_outputs_2_PENABLE <= io_input_PENABLE;
  io_outputs_2_PSEL(0) <= pkg_extract(io_input_PSEL,2);
  io_outputs_2_PWRITE <= io_input_PWRITE;
  io_outputs_2_PWDATA <= io_input_PWDATA;
  zz_selIndex <= pkg_extract(io_input_PSEL,1);
  zz_selIndex_1 <= pkg_extract(io_input_PSEL,2);
  io_input_PREADY <= zz_io_input_PREADY;
  io_input_PRDATA <= zz_io_input_PRDATA;
  io_input_PSLVERROR <= zz_io_input_PSLVERROR;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      selIndex <= unsigned(pkg_cat(pkg_toStdLogicVector(zz_selIndex_1),pkg_toStdLogicVector(zz_selIndex)));
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity Muraxy is
  port(
    io_asyncReset : in std_logic;
    io_mainClk : in std_logic;
    io_gpioA_read : in std_logic_vector(31 downto 0);
    io_gpioA_write : out std_logic_vector(31 downto 0);
    io_gpioA_writeEnable : out std_logic_vector(31 downto 0);
    io_uart_txd : out std_logic;
    io_uart_rxd : in std_logic
  );
end Muraxy;

architecture arch of Muraxy is
  signal axi_gpioACtrl_io_apb_PADDR : unsigned(3 downto 0);
  signal axi_uartCtrl_io_apb_PADDR : unsigned(4 downto 0);
  signal axi_timer_io_apb_PADDR : unsigned(7 downto 0);
  signal axi_core_cpu_dBus_cmd_ready : std_logic;
  signal axi_core_cpu_dBus_rsp_payload_last : std_logic;
  signal axi_core_cpu_dBus_rsp_payload_error : std_logic;
  signal axi_core_cpu_debug_bus_cmd_payload_address : unsigned(7 downto 0);
  signal axi_core_cpu_iBus_rsp_payload_error : std_logic;
  signal streamFork_3_io_input_valid : std_logic;
  signal streamFork_3_io_outputs_0_ready : std_logic;
  signal streamFork_3_io_outputs_1_ready : std_logic;
  signal dbus_axi_decoder_io_input_r_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr : unsigned(14 downto 0);
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_arw_payload_addr : unsigned(14 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_arw_payload_addr : unsigned(19 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_ready : std_logic;
  signal io_asyncReset_buffercc_io_dataOut : std_logic;
  signal axi_ram_io_axi_arw_ready : std_logic;
  signal axi_ram_io_axi_w_ready : std_logic;
  signal axi_ram_io_axi_b_valid : std_logic;
  signal axi_ram_io_axi_b_payload_id : unsigned(3 downto 0);
  signal axi_ram_io_axi_b_payload_resp : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_r_valid : std_logic;
  signal axi_ram_io_axi_r_payload_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_r_payload_id : unsigned(3 downto 0);
  signal axi_ram_io_axi_r_payload_resp : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_r_payload_last : std_logic;
  signal axi_apbBridge_io_axi_arw_ready : std_logic;
  signal axi_apbBridge_io_axi_w_ready : std_logic;
  signal axi_apbBridge_io_axi_b_valid : std_logic;
  signal axi_apbBridge_io_axi_b_payload_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_b_payload_resp : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_r_valid : std_logic;
  signal axi_apbBridge_io_axi_r_payload_data : std_logic_vector(31 downto 0);
  signal axi_apbBridge_io_axi_r_payload_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_r_payload_resp : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_r_payload_last : std_logic;
  signal axi_apbBridge_io_apb_PADDR : unsigned(19 downto 0);
  signal axi_apbBridge_io_apb_PSEL : std_logic_vector(0 downto 0);
  signal axi_apbBridge_io_apb_PENABLE : std_logic;
  signal axi_apbBridge_io_apb_PWRITE : std_logic;
  signal axi_apbBridge_io_apb_PWDATA : std_logic_vector(31 downto 0);
  signal axi_gpioACtrl_io_apb_PREADY : std_logic;
  signal axi_gpioACtrl_io_apb_PRDATA : std_logic_vector(31 downto 0);
  signal axi_gpioACtrl_io_apb_PSLVERROR : std_logic;
  signal axi_gpioACtrl_io_gpio_write : std_logic_vector(31 downto 0);
  signal axi_gpioACtrl_io_gpio_writeEnable : std_logic_vector(31 downto 0);
  signal axi_gpioACtrl_io_value : std_logic_vector(31 downto 0);
  signal axi_uartCtrl_io_apb_PREADY : std_logic;
  signal axi_uartCtrl_io_apb_PRDATA : std_logic_vector(31 downto 0);
  signal axi_uartCtrl_io_uart_txd : std_logic;
  signal axi_uartCtrl_io_interrupt : std_logic;
  signal axi_timer_io_apb_PREADY : std_logic;
  signal axi_timer_io_apb_PRDATA : std_logic_vector(31 downto 0);
  signal axi_timer_io_apb_PSLVERROR : std_logic;
  signal axi_timer_io_interrupt : std_logic;
  signal axi_core_cpu_dBus_cmd_valid : std_logic;
  signal axi_core_cpu_dBus_cmd_payload_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_payload_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_payload_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_payload_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_payload_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_payload_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_payload_last : std_logic;
  signal axi_core_cpu_debug_bus_cmd_ready : std_logic;
  signal axi_core_cpu_debug_bus_rsp_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_debug_resetOut : std_logic;
  signal axi_core_cpu_iBus_cmd_valid : std_logic;
  signal axi_core_cpu_iBus_cmd_payload_address : unsigned(31 downto 0);
  signal axi_core_cpu_iBus_cmd_payload_size : unsigned(2 downto 0);
  signal streamFork_3_io_input_ready : std_logic;
  signal streamFork_3_io_outputs_0_valid : std_logic;
  signal streamFork_3_io_outputs_0_payload_wr : std_logic;
  signal streamFork_3_io_outputs_0_payload_uncached : std_logic;
  signal streamFork_3_io_outputs_0_payload_address : unsigned(31 downto 0);
  signal streamFork_3_io_outputs_0_payload_data : std_logic_vector(31 downto 0);
  signal streamFork_3_io_outputs_0_payload_mask : std_logic_vector(3 downto 0);
  signal streamFork_3_io_outputs_0_payload_size : unsigned(2 downto 0);
  signal streamFork_3_io_outputs_0_payload_last : std_logic;
  signal streamFork_3_io_outputs_1_valid : std_logic;
  signal streamFork_3_io_outputs_1_payload_wr : std_logic;
  signal streamFork_3_io_outputs_1_payload_uncached : std_logic;
  signal streamFork_3_io_outputs_1_payload_address : unsigned(31 downto 0);
  signal streamFork_3_io_outputs_1_payload_data : std_logic_vector(31 downto 0);
  signal streamFork_3_io_outputs_1_payload_mask : std_logic_vector(3 downto 0);
  signal streamFork_3_io_outputs_1_payload_size : unsigned(2 downto 0);
  signal streamFork_3_io_outputs_1_payload_last : std_logic;
  signal bSCANE2_1_CAPTURE : std_logic;
  signal bSCANE2_1_DRCK : std_logic;
  signal bSCANE2_1_RESET : std_logic;
  signal bSCANE2_1_RUNTEST : std_logic;
  signal bSCANE2_1_SEL : std_logic;
  signal bSCANE2_1_SHIFT : std_logic;
  signal bSCANE2_1_TCK : std_logic;
  signal bSCANE2_1_TDI : std_logic;
  signal bSCANE2_1_TMS : std_logic;
  signal bSCANE2_1_UPDATE : std_logic;
  signal jtagBridgeNoTap_1_io_ctrl_tdo : std_logic;
  signal jtagBridgeNoTap_1_io_remote_cmd_valid : std_logic;
  signal jtagBridgeNoTap_1_io_remote_cmd_payload_last : std_logic;
  signal jtagBridgeNoTap_1_io_remote_cmd_payload_fragment : std_logic_vector(0 downto 0);
  signal jtagBridgeNoTap_1_io_remote_rsp_ready : std_logic;
  signal systemDebugger_1_io_remote_cmd_ready : std_logic;
  signal systemDebugger_1_io_remote_rsp_valid : std_logic;
  signal systemDebugger_1_io_remote_rsp_payload_error : std_logic;
  signal systemDebugger_1_io_remote_rsp_payload_data : std_logic_vector(31 downto 0);
  signal systemDebugger_1_io_mem_cmd_valid : std_logic;
  signal systemDebugger_1_io_mem_cmd_payload_address : unsigned(31 downto 0);
  signal systemDebugger_1_io_mem_cmd_payload_data : std_logic_vector(31 downto 0);
  signal systemDebugger_1_io_mem_cmd_payload_wr : std_logic;
  signal systemDebugger_1_io_mem_cmd_payload_size : unsigned(1 downto 0);
  signal axi4ReadOnlyDecoder_1_io_input_ar_ready : std_logic;
  signal axi4ReadOnlyDecoder_1_io_input_r_valid : std_logic;
  signal axi4ReadOnlyDecoder_1_io_input_r_payload_data : std_logic_vector(31 downto 0);
  signal axi4ReadOnlyDecoder_1_io_input_r_payload_resp : std_logic_vector(1 downto 0);
  signal axi4ReadOnlyDecoder_1_io_input_r_payload_last : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_valid : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_addr : unsigned(31 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_len : unsigned(7 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_burst : std_logic_vector(1 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_cache : std_logic_vector(3 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_prot : std_logic_vector(2 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_r_ready : std_logic;
  signal dbus_axi_decoder_io_input_arw_ready : std_logic;
  signal dbus_axi_decoder_io_input_w_ready : std_logic;
  signal dbus_axi_decoder_io_input_b_valid : std_logic;
  signal dbus_axi_decoder_io_input_b_payload_resp : std_logic_vector(1 downto 0);
  signal dbus_axi_decoder_io_input_r_valid : std_logic;
  signal dbus_axi_decoder_io_input_r_payload_data : std_logic_vector(31 downto 0);
  signal dbus_axi_decoder_io_input_r_payload_resp : std_logic_vector(1 downto 0);
  signal dbus_axi_decoder_io_input_r_payload_last : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_valid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_payload_addr : unsigned(31 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_payload_len : unsigned(7 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_payload_size : unsigned(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_payload_cache : std_logic_vector(3 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_payload_prot : std_logic_vector(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_payload_write : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_w_valid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_w_payload_data : std_logic_vector(31 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_w_payload_strb : std_logic_vector(3 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_w_payload_last : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_b_ready : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_r_ready : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_valid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_payload_addr : unsigned(31 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_payload_len : unsigned(7 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_payload_size : unsigned(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_payload_cache : std_logic_vector(3 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_payload_prot : std_logic_vector(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_payload_write : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_w_valid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_w_payload_data : std_logic_vector(31 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_w_payload_strb : std_logic_vector(3 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_w_payload_last : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_b_ready : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_r_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_readInputs_0_ar_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_readInputs_0_r_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_id : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_resp : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_last : std_logic;
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_arw_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_w_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_b_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_b_payload_id : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_b_payload_resp : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_r_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_id : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_resp : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_last : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_payload_addr : unsigned(14 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_payload_id : unsigned(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_payload_len : unsigned(7 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_payload_size : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_payload_burst : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_payload_write : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_payload_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_payload_strb : std_logic_vector(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_payload_last : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_b_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_r_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_arw_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_w_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_valid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_payload_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_payload_resp : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_valid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_data : std_logic_vector(31 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_resp : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_last : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_valid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_payload_addr : unsigned(19 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_payload_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_payload_len : unsigned(7 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_payload_size : unsigned(2 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_payload_burst : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_payload_write : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_valid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_payload_data : std_logic_vector(31 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_w_payload_strb : std_logic_vector(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_w_payload_last : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_b_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_r_ready : std_logic;
  signal io_apb_decoder_io_input_PREADY : std_logic;
  signal io_apb_decoder_io_input_PRDATA : std_logic_vector(31 downto 0);
  signal io_apb_decoder_io_input_PSLVERROR : std_logic;
  signal io_apb_decoder_io_output_PADDR : unsigned(19 downto 0);
  signal io_apb_decoder_io_output_PSEL : std_logic_vector(2 downto 0);
  signal io_apb_decoder_io_output_PENABLE : std_logic;
  signal io_apb_decoder_io_output_PWRITE : std_logic;
  signal io_apb_decoder_io_output_PWDATA : std_logic_vector(31 downto 0);
  signal apb3Router_1_io_input_PREADY : std_logic;
  signal apb3Router_1_io_input_PRDATA : std_logic_vector(31 downto 0);
  signal apb3Router_1_io_input_PSLVERROR : std_logic;
  signal apb3Router_1_io_outputs_0_PADDR : unsigned(19 downto 0);
  signal apb3Router_1_io_outputs_0_PSEL : std_logic_vector(0 downto 0);
  signal apb3Router_1_io_outputs_0_PENABLE : std_logic;
  signal apb3Router_1_io_outputs_0_PWRITE : std_logic;
  signal apb3Router_1_io_outputs_0_PWDATA : std_logic_vector(31 downto 0);
  signal apb3Router_1_io_outputs_1_PADDR : unsigned(19 downto 0);
  signal apb3Router_1_io_outputs_1_PSEL : std_logic_vector(0 downto 0);
  signal apb3Router_1_io_outputs_1_PENABLE : std_logic;
  signal apb3Router_1_io_outputs_1_PWRITE : std_logic;
  signal apb3Router_1_io_outputs_1_PWDATA : std_logic_vector(31 downto 0);
  signal apb3Router_1_io_outputs_2_PADDR : unsigned(19 downto 0);
  signal apb3Router_1_io_outputs_2_PSEL : std_logic_vector(0 downto 0);
  signal apb3Router_1_io_outputs_2_PENABLE : std_logic;
  signal apb3Router_1_io_outputs_2_PWRITE : std_logic;
  signal apb3Router_1_io_outputs_2_PWDATA : std_logic_vector(31 downto 0);

  component BSCANE2 is
    generic( 
      DISABLE_JTAG : string ;
      JTAG_CHAIN : integer  
    );
    port( 
      CAPTURE : out std_logic;
      DRCK : out std_logic;
      RESET : out std_logic;
      RUNTEST : out std_logic;
      SEL : out std_logic;
      SHIFT : out std_logic;
      TCK : out std_logic;
      TDI : out std_logic;
      TMS : out std_logic;
      UPDATE : out std_logic;
      TDO : in std_logic 
    );
  end component;
  

  signal resetCtrl_systemResetUnbuffered : std_logic;
  signal resetCtrl_systemResetCounter : unsigned(5 downto 0) := pkg_unsigned("000000");
  signal zz_when_Muraxy_l198 : unsigned(5 downto 0);
  signal when_Muraxy_l198 : std_logic;
  signal when_Muraxy_l202 : std_logic;
  signal resetCtrl_systemReset : std_logic;
  signal resetCtrl_axiReset : std_logic;
  signal dbus_axi_arw_valid : std_logic;
  signal dbus_axi_arw_ready : std_logic;
  signal dbus_axi_arw_payload_addr : unsigned(31 downto 0);
  signal dbus_axi_arw_payload_len : unsigned(7 downto 0);
  signal dbus_axi_arw_payload_size : unsigned(2 downto 0);
  signal dbus_axi_arw_payload_cache : std_logic_vector(3 downto 0);
  signal dbus_axi_arw_payload_prot : std_logic_vector(2 downto 0);
  signal dbus_axi_arw_payload_write : std_logic;
  signal dbus_axi_w_valid : std_logic;
  signal dbus_axi_w_ready : std_logic;
  signal dbus_axi_w_payload_data : std_logic_vector(31 downto 0);
  signal dbus_axi_w_payload_strb : std_logic_vector(3 downto 0);
  signal dbus_axi_w_payload_last : std_logic;
  signal dbus_axi_b_valid : std_logic;
  signal dbus_axi_b_ready : std_logic;
  signal dbus_axi_b_payload_resp : std_logic_vector(1 downto 0);
  signal dbus_axi_r_valid : std_logic;
  signal dbus_axi_r_ready : std_logic;
  signal dbus_axi_r_payload_data : std_logic_vector(31 downto 0);
  signal dbus_axi_r_payload_resp : std_logic_vector(1 downto 0);
  signal dbus_axi_r_payload_last : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_valid : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_ready : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_payload_last : std_logic;
  signal axi_core_cpu_dBus_cmd_rValid : std_logic;
  signal axi_core_cpu_dBus_cmd_rData_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_rData_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_rData_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_rData_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_rData_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_rData_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_rData_last : std_logic;
  signal when_Stream_l342 : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_valid : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_ready : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_last : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_rValid : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_rData_last : std_logic;
  signal when_Stream_l342_1 : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_valid : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_last : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_wr : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_uncached : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_address : unsigned(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_data : std_logic_vector(31 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_mask : std_logic_vector(3 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_size : unsigned(2 downto 0);
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_last : std_logic;
  signal axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_fire : std_logic;
  signal when_Utils_l594 : std_logic;
  signal dbus_axi_b_fire : std_logic;
  signal zz_when_Utils_l622 : std_logic;
  signal zz_when_Utils_l622_1 : std_logic;
  signal zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready : unsigned(2 downto 0);
  signal zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_1 : unsigned(2 downto 0);
  signal when_Utils_l622 : std_logic;
  signal when_Utils_l624 : std_logic;
  signal zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_2 : std_logic;
  signal streamFork_3_io_outputs_0_fire : std_logic;
  signal zz_1 : std_logic;
  signal streamFork_3_io_outputs_0_thrown_valid : std_logic;
  signal streamFork_3_io_outputs_0_thrown_ready : std_logic;
  signal streamFork_3_io_outputs_0_thrown_payload_wr : std_logic;
  signal streamFork_3_io_outputs_0_thrown_payload_uncached : std_logic;
  signal streamFork_3_io_outputs_0_thrown_payload_address : unsigned(31 downto 0);
  signal streamFork_3_io_outputs_0_thrown_payload_data : std_logic_vector(31 downto 0);
  signal streamFork_3_io_outputs_0_thrown_payload_mask : std_logic_vector(3 downto 0);
  signal streamFork_3_io_outputs_0_thrown_payload_size : unsigned(2 downto 0);
  signal streamFork_3_io_outputs_0_thrown_payload_last : std_logic;
  signal when_Stream_l408 : std_logic;
  signal streamFork_3_io_outputs_1_thrown_valid : std_logic;
  signal streamFork_3_io_outputs_1_thrown_ready : std_logic;
  signal streamFork_3_io_outputs_1_thrown_payload_wr : std_logic;
  signal streamFork_3_io_outputs_1_thrown_payload_uncached : std_logic;
  signal streamFork_3_io_outputs_1_thrown_payload_address : unsigned(31 downto 0);
  signal streamFork_3_io_outputs_1_thrown_payload_data : std_logic_vector(31 downto 0);
  signal streamFork_3_io_outputs_1_thrown_payload_mask : std_logic_vector(3 downto 0);
  signal streamFork_3_io_outputs_1_thrown_payload_size : unsigned(2 downto 0);
  signal streamFork_3_io_outputs_1_thrown_payload_last : std_logic;
  signal axi_core_cpu_debug_resetOut_regNext : std_logic;
  signal axi_core_cpu_debug_bus_cmd_fire : std_logic;
  signal axi_core_cpu_debug_bus_cmd_fire_regNext : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_valid : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_ready : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_addr : unsigned(31 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_len : unsigned(7 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_burst : std_logic_vector(1 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_cache : std_logic_vector(3 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_prot : std_logic_vector(2 downto 0);
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_rValid : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_fire : std_logic;
  signal axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_fire_1 : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_valid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_ready : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_addr : unsigned(31 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_len : unsigned(7 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_size : unsigned(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_cache : std_logic_vector(3 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_prot : std_logic_vector(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_write : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_rValid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_fire : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_fire_1 : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_valid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_ready : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_addr : unsigned(31 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_len : unsigned(7 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_size : unsigned(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_cache : std_logic_vector(3 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_prot : std_logic_vector(2 downto 0);
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_write : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_rValid : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_fire : std_logic;
  signal dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_fire_1 : std_logic;
  signal dbus_axi_decoder_io_input_r_m2sPipe_valid : std_logic;
  signal dbus_axi_decoder_io_input_r_m2sPipe_ready : std_logic;
  signal dbus_axi_decoder_io_input_r_m2sPipe_payload_data : std_logic_vector(31 downto 0);
  signal dbus_axi_decoder_io_input_r_m2sPipe_payload_resp : std_logic_vector(1 downto 0);
  signal dbus_axi_decoder_io_input_r_m2sPipe_payload_last : std_logic;
  signal dbus_axi_decoder_io_input_r_rValid : std_logic;
  signal dbus_axi_decoder_io_input_r_rData_data : std_logic_vector(31 downto 0);
  signal dbus_axi_decoder_io_input_r_rData_resp : std_logic_vector(1 downto 0);
  signal dbus_axi_decoder_io_input_r_rData_last : std_logic;
  signal when_Stream_l342_2 : std_logic;
  signal zz_io_readInputs_0_ar_payload_id : unsigned(2 downto 0);
  signal zz_io_sharedInputs_0_arw_payload_id : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_addr : unsigned(14 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_id : unsigned(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_len : unsigned(7 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_size : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_burst : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_write : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_rValid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_halfPipe_fire : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_arw_rData_addr : unsigned(14 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_rData_id : unsigned(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_rData_len : unsigned(7 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_rData_size : unsigned(2 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_rData_burst : std_logic_vector(1 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_arw_rData_write : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_strb : std_logic_vector(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_last : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_rValid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_rData_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_rData_strb : std_logic_vector(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_rData_last : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_valid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_ready : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_strb : std_logic_vector(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_last : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rValid : std_logic;
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_data : std_logic_vector(31 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_strb : std_logic_vector(3 downto 0);
  signal axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_last : std_logic;
  signal when_Stream_l342_3 : std_logic;
  signal zz_io_sharedInputs_0_arw_payload_id_1 : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_valid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_addr : unsigned(19 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_len : unsigned(7 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_size : unsigned(2 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_burst : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_write : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rValid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_fire : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rData_addr : unsigned(19 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rData_id : unsigned(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rData_len : unsigned(7 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rData_size : unsigned(2 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rData_burst : std_logic_vector(1 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_arw_rData_write : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_valid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_ready : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_data : std_logic_vector(31 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_strb : std_logic_vector(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_last : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_rValid : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_fire : std_logic;
  signal axi_apbBridge_io_axi_arbiter_io_output_w_rData_data : std_logic_vector(31 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_w_rData_strb : std_logic_vector(3 downto 0);
  signal axi_apbBridge_io_axi_arbiter_io_output_w_rData_last : std_logic;
begin
  io_asyncReset_buffercc : entity work.BufferCC_3
    port map ( 
      io_dataIn => io_asyncReset,
      io_dataOut => io_asyncReset_buffercc_io_dataOut,
      io_mainClk => io_mainClk 
    );
  axi_ram : entity work.Axi4SharedOnChipRam
    port map ( 
      io_axi_arw_valid => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_valid,
      io_axi_arw_ready => axi_ram_io_axi_arw_ready,
      io_axi_arw_payload_addr => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_addr,
      io_axi_arw_payload_id => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_id,
      io_axi_arw_payload_len => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_len,
      io_axi_arw_payload_size => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_size,
      io_axi_arw_payload_burst => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_burst,
      io_axi_arw_payload_write => axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_write,
      io_axi_w_valid => axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_valid,
      io_axi_w_ready => axi_ram_io_axi_w_ready,
      io_axi_w_payload_data => axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_data,
      io_axi_w_payload_strb => axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_strb,
      io_axi_w_payload_last => axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_last,
      io_axi_b_valid => axi_ram_io_axi_b_valid,
      io_axi_b_ready => axi_ram_io_axi_arbiter_io_output_b_ready,
      io_axi_b_payload_id => axi_ram_io_axi_b_payload_id,
      io_axi_b_payload_resp => axi_ram_io_axi_b_payload_resp,
      io_axi_r_valid => axi_ram_io_axi_r_valid,
      io_axi_r_ready => axi_ram_io_axi_arbiter_io_output_r_ready,
      io_axi_r_payload_data => axi_ram_io_axi_r_payload_data,
      io_axi_r_payload_id => axi_ram_io_axi_r_payload_id,
      io_axi_r_payload_resp => axi_ram_io_axi_r_payload_resp,
      io_axi_r_payload_last => axi_ram_io_axi_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_apbBridge : entity work.Axi4SharedToApb3Bridge
    port map ( 
      io_axi_arw_valid => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_valid,
      io_axi_arw_ready => axi_apbBridge_io_axi_arw_ready,
      io_axi_arw_payload_addr => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_addr,
      io_axi_arw_payload_id => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_id,
      io_axi_arw_payload_len => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_len,
      io_axi_arw_payload_size => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_size,
      io_axi_arw_payload_burst => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_burst,
      io_axi_arw_payload_write => axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_write,
      io_axi_w_valid => axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_valid,
      io_axi_w_ready => axi_apbBridge_io_axi_w_ready,
      io_axi_w_payload_data => axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_data,
      io_axi_w_payload_strb => axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_strb,
      io_axi_w_payload_last => axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_last,
      io_axi_b_valid => axi_apbBridge_io_axi_b_valid,
      io_axi_b_ready => axi_apbBridge_io_axi_arbiter_io_output_b_ready,
      io_axi_b_payload_id => axi_apbBridge_io_axi_b_payload_id,
      io_axi_b_payload_resp => axi_apbBridge_io_axi_b_payload_resp,
      io_axi_r_valid => axi_apbBridge_io_axi_r_valid,
      io_axi_r_ready => axi_apbBridge_io_axi_arbiter_io_output_r_ready,
      io_axi_r_payload_data => axi_apbBridge_io_axi_r_payload_data,
      io_axi_r_payload_id => axi_apbBridge_io_axi_r_payload_id,
      io_axi_r_payload_resp => axi_apbBridge_io_axi_r_payload_resp,
      io_axi_r_payload_last => axi_apbBridge_io_axi_r_payload_last,
      io_apb_PADDR => axi_apbBridge_io_apb_PADDR,
      io_apb_PSEL => axi_apbBridge_io_apb_PSEL,
      io_apb_PENABLE => axi_apbBridge_io_apb_PENABLE,
      io_apb_PREADY => io_apb_decoder_io_input_PREADY,
      io_apb_PWRITE => axi_apbBridge_io_apb_PWRITE,
      io_apb_PWDATA => axi_apbBridge_io_apb_PWDATA,
      io_apb_PRDATA => io_apb_decoder_io_input_PRDATA,
      io_apb_PSLVERROR => io_apb_decoder_io_input_PSLVERROR,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_gpioACtrl : entity work.Apb3Gpio
    port map ( 
      io_apb_PADDR => axi_gpioACtrl_io_apb_PADDR,
      io_apb_PSEL => apb3Router_1_io_outputs_0_PSEL,
      io_apb_PENABLE => apb3Router_1_io_outputs_0_PENABLE,
      io_apb_PREADY => axi_gpioACtrl_io_apb_PREADY,
      io_apb_PWRITE => apb3Router_1_io_outputs_0_PWRITE,
      io_apb_PWDATA => apb3Router_1_io_outputs_0_PWDATA,
      io_apb_PRDATA => axi_gpioACtrl_io_apb_PRDATA,
      io_apb_PSLVERROR => axi_gpioACtrl_io_apb_PSLVERROR,
      io_gpio_read => io_gpioA_read,
      io_gpio_write => axi_gpioACtrl_io_gpio_write,
      io_gpio_writeEnable => axi_gpioACtrl_io_gpio_writeEnable,
      io_value => axi_gpioACtrl_io_value,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_uartCtrl : entity work.Apb3UartCtrl
    port map ( 
      io_apb_PADDR => axi_uartCtrl_io_apb_PADDR,
      io_apb_PSEL => apb3Router_1_io_outputs_1_PSEL,
      io_apb_PENABLE => apb3Router_1_io_outputs_1_PENABLE,
      io_apb_PREADY => axi_uartCtrl_io_apb_PREADY,
      io_apb_PWRITE => apb3Router_1_io_outputs_1_PWRITE,
      io_apb_PWDATA => apb3Router_1_io_outputs_1_PWDATA,
      io_apb_PRDATA => axi_uartCtrl_io_apb_PRDATA,
      io_uart_txd => axi_uartCtrl_io_uart_txd,
      io_uart_rxd => io_uart_rxd,
      io_interrupt => axi_uartCtrl_io_interrupt,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_timer : entity work.MuraxApb3Timer
    port map ( 
      io_apb_PADDR => axi_timer_io_apb_PADDR,
      io_apb_PSEL => apb3Router_1_io_outputs_2_PSEL,
      io_apb_PENABLE => apb3Router_1_io_outputs_2_PENABLE,
      io_apb_PREADY => axi_timer_io_apb_PREADY,
      io_apb_PWRITE => apb3Router_1_io_outputs_2_PWRITE,
      io_apb_PWDATA => apb3Router_1_io_outputs_2_PWDATA,
      io_apb_PRDATA => axi_timer_io_apb_PRDATA,
      io_apb_PSLVERROR => axi_timer_io_apb_PSLVERROR,
      io_interrupt => axi_timer_io_interrupt,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_core_cpu : entity work.VexRiscv
    port map ( 
      dBus_cmd_valid => axi_core_cpu_dBus_cmd_valid,
      dBus_cmd_ready => axi_core_cpu_dBus_cmd_ready,
      dBus_cmd_payload_wr => axi_core_cpu_dBus_cmd_payload_wr,
      dBus_cmd_payload_uncached => axi_core_cpu_dBus_cmd_payload_uncached,
      dBus_cmd_payload_address => axi_core_cpu_dBus_cmd_payload_address,
      dBus_cmd_payload_data => axi_core_cpu_dBus_cmd_payload_data,
      dBus_cmd_payload_mask => axi_core_cpu_dBus_cmd_payload_mask,
      dBus_cmd_payload_size => axi_core_cpu_dBus_cmd_payload_size,
      dBus_cmd_payload_last => axi_core_cpu_dBus_cmd_payload_last,
      dBus_rsp_valid => dbus_axi_r_valid,
      dBus_rsp_payload_last => axi_core_cpu_dBus_rsp_payload_last,
      dBus_rsp_payload_data => dbus_axi_r_payload_data,
      dBus_rsp_payload_error => axi_core_cpu_dBus_rsp_payload_error,
      timerInterrupt => axi_timer_io_interrupt,
      externalInterrupt => pkg_toStdLogic(false),
      softwareInterrupt => pkg_toStdLogic(false),
      debug_bus_cmd_valid => systemDebugger_1_io_mem_cmd_valid,
      debug_bus_cmd_ready => axi_core_cpu_debug_bus_cmd_ready,
      debug_bus_cmd_payload_wr => systemDebugger_1_io_mem_cmd_payload_wr,
      debug_bus_cmd_payload_address => axi_core_cpu_debug_bus_cmd_payload_address,
      debug_bus_cmd_payload_data => systemDebugger_1_io_mem_cmd_payload_data,
      debug_bus_rsp_data => axi_core_cpu_debug_bus_rsp_data,
      debug_resetOut => axi_core_cpu_debug_resetOut,
      iBus_cmd_valid => axi_core_cpu_iBus_cmd_valid,
      iBus_cmd_ready => axi4ReadOnlyDecoder_1_io_input_ar_ready,
      iBus_cmd_payload_address => axi_core_cpu_iBus_cmd_payload_address,
      iBus_cmd_payload_size => axi_core_cpu_iBus_cmd_payload_size,
      iBus_rsp_valid => axi4ReadOnlyDecoder_1_io_input_r_valid,
      iBus_rsp_payload_data => axi4ReadOnlyDecoder_1_io_input_r_payload_data,
      iBus_rsp_payload_error => axi_core_cpu_iBus_rsp_payload_error,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset,
      resetCtrl_systemReset => resetCtrl_systemReset 
    );
  streamFork_3 : entity work.StreamFork_2
    port map ( 
      io_input_valid => streamFork_3_io_input_valid,
      io_input_ready => streamFork_3_io_input_ready,
      io_input_payload_wr => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_wr,
      io_input_payload_uncached => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_uncached,
      io_input_payload_address => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_address,
      io_input_payload_data => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_data,
      io_input_payload_mask => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_mask,
      io_input_payload_size => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_size,
      io_input_payload_last => axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_last,
      io_outputs_0_valid => streamFork_3_io_outputs_0_valid,
      io_outputs_0_ready => streamFork_3_io_outputs_0_ready,
      io_outputs_0_payload_wr => streamFork_3_io_outputs_0_payload_wr,
      io_outputs_0_payload_uncached => streamFork_3_io_outputs_0_payload_uncached,
      io_outputs_0_payload_address => streamFork_3_io_outputs_0_payload_address,
      io_outputs_0_payload_data => streamFork_3_io_outputs_0_payload_data,
      io_outputs_0_payload_mask => streamFork_3_io_outputs_0_payload_mask,
      io_outputs_0_payload_size => streamFork_3_io_outputs_0_payload_size,
      io_outputs_0_payload_last => streamFork_3_io_outputs_0_payload_last,
      io_outputs_1_valid => streamFork_3_io_outputs_1_valid,
      io_outputs_1_ready => streamFork_3_io_outputs_1_ready,
      io_outputs_1_payload_wr => streamFork_3_io_outputs_1_payload_wr,
      io_outputs_1_payload_uncached => streamFork_3_io_outputs_1_payload_uncached,
      io_outputs_1_payload_address => streamFork_3_io_outputs_1_payload_address,
      io_outputs_1_payload_data => streamFork_3_io_outputs_1_payload_data,
      io_outputs_1_payload_mask => streamFork_3_io_outputs_1_payload_mask,
      io_outputs_1_payload_size => streamFork_3_io_outputs_1_payload_size,
      io_outputs_1_payload_last => streamFork_3_io_outputs_1_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  bSCANE2_1 : BSCANE2
    generic map( 
      DISABLE_JTAG => "FALSE",
      JTAG_CHAIN => 2 
    )
    port map ( 
      CAPTURE => bSCANE2_1_CAPTURE,
      DRCK => bSCANE2_1_DRCK,
      RESET => bSCANE2_1_RESET,
      RUNTEST => bSCANE2_1_RUNTEST,
      SEL => bSCANE2_1_SEL,
      SHIFT => bSCANE2_1_SHIFT,
      TCK => bSCANE2_1_TCK,
      TDI => bSCANE2_1_TDI,
      TMS => bSCANE2_1_TMS,
      UPDATE => bSCANE2_1_UPDATE,
      TDO => jtagBridgeNoTap_1_io_ctrl_tdo 
    );
  jtagBridgeNoTap_1 : entity work.JtagBridgeNoTap
    port map ( 
      io_ctrl_tdi => bSCANE2_1_TDI,
      io_ctrl_enable => bSCANE2_1_SEL,
      io_ctrl_capture => bSCANE2_1_CAPTURE,
      io_ctrl_shift => bSCANE2_1_SHIFT,
      io_ctrl_update => bSCANE2_1_UPDATE,
      io_ctrl_reset => bSCANE2_1_RESET,
      io_ctrl_tdo => jtagBridgeNoTap_1_io_ctrl_tdo,
      io_remote_cmd_valid => jtagBridgeNoTap_1_io_remote_cmd_valid,
      io_remote_cmd_ready => systemDebugger_1_io_remote_cmd_ready,
      io_remote_cmd_payload_last => jtagBridgeNoTap_1_io_remote_cmd_payload_last,
      io_remote_cmd_payload_fragment => jtagBridgeNoTap_1_io_remote_cmd_payload_fragment,
      io_remote_rsp_valid => systemDebugger_1_io_remote_rsp_valid,
      io_remote_rsp_ready => jtagBridgeNoTap_1_io_remote_rsp_ready,
      io_remote_rsp_payload_error => systemDebugger_1_io_remote_rsp_payload_error,
      io_remote_rsp_payload_data => systemDebugger_1_io_remote_rsp_payload_data,
      io_mainClk => io_mainClk,
      resetCtrl_systemReset => resetCtrl_systemReset,
      TCK => bSCANE2_1_TCK 
    );
  systemDebugger_1 : entity work.SystemDebugger
    port map ( 
      io_remote_cmd_valid => jtagBridgeNoTap_1_io_remote_cmd_valid,
      io_remote_cmd_ready => systemDebugger_1_io_remote_cmd_ready,
      io_remote_cmd_payload_last => jtagBridgeNoTap_1_io_remote_cmd_payload_last,
      io_remote_cmd_payload_fragment => jtagBridgeNoTap_1_io_remote_cmd_payload_fragment,
      io_remote_rsp_valid => systemDebugger_1_io_remote_rsp_valid,
      io_remote_rsp_ready => jtagBridgeNoTap_1_io_remote_rsp_ready,
      io_remote_rsp_payload_error => systemDebugger_1_io_remote_rsp_payload_error,
      io_remote_rsp_payload_data => systemDebugger_1_io_remote_rsp_payload_data,
      io_mem_cmd_valid => systemDebugger_1_io_mem_cmd_valid,
      io_mem_cmd_ready => axi_core_cpu_debug_bus_cmd_ready,
      io_mem_cmd_payload_address => systemDebugger_1_io_mem_cmd_payload_address,
      io_mem_cmd_payload_data => systemDebugger_1_io_mem_cmd_payload_data,
      io_mem_cmd_payload_wr => systemDebugger_1_io_mem_cmd_payload_wr,
      io_mem_cmd_payload_size => systemDebugger_1_io_mem_cmd_payload_size,
      io_mem_rsp_valid => axi_core_cpu_debug_bus_cmd_fire_regNext,
      io_mem_rsp_payload => axi_core_cpu_debug_bus_rsp_data,
      io_mainClk => io_mainClk,
      resetCtrl_systemReset => resetCtrl_systemReset 
    );
  axi4ReadOnlyDecoder_1 : entity work.Axi4ReadOnlyDecoder
    port map ( 
      io_input_ar_valid => axi_core_cpu_iBus_cmd_valid,
      io_input_ar_ready => axi4ReadOnlyDecoder_1_io_input_ar_ready,
      io_input_ar_payload_addr => axi_core_cpu_iBus_cmd_payload_address,
      io_input_ar_payload_len => pkg_unsigned("00000111"),
      io_input_ar_payload_burst => pkg_stdLogicVector("01"),
      io_input_ar_payload_cache => pkg_stdLogicVector("1111"),
      io_input_ar_payload_prot => pkg_stdLogicVector("110"),
      io_input_r_valid => axi4ReadOnlyDecoder_1_io_input_r_valid,
      io_input_r_ready => pkg_toStdLogic(true),
      io_input_r_payload_data => axi4ReadOnlyDecoder_1_io_input_r_payload_data,
      io_input_r_payload_resp => axi4ReadOnlyDecoder_1_io_input_r_payload_resp,
      io_input_r_payload_last => axi4ReadOnlyDecoder_1_io_input_r_payload_last,
      io_outputs_0_ar_valid => axi4ReadOnlyDecoder_1_io_outputs_0_ar_valid,
      io_outputs_0_ar_ready => axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_fire_1,
      io_outputs_0_ar_payload_addr => axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_addr,
      io_outputs_0_ar_payload_len => axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_len,
      io_outputs_0_ar_payload_burst => axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_burst,
      io_outputs_0_ar_payload_cache => axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_cache,
      io_outputs_0_ar_payload_prot => axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_prot,
      io_outputs_0_r_valid => axi_ram_io_axi_arbiter_io_readInputs_0_r_valid,
      io_outputs_0_r_ready => axi4ReadOnlyDecoder_1_io_outputs_0_r_ready,
      io_outputs_0_r_payload_data => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_data,
      io_outputs_0_r_payload_resp => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_resp,
      io_outputs_0_r_payload_last => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  dbus_axi_decoder : entity work.Axi4SharedDecoder
    port map ( 
      io_input_arw_valid => dbus_axi_arw_valid,
      io_input_arw_ready => dbus_axi_decoder_io_input_arw_ready,
      io_input_arw_payload_addr => dbus_axi_arw_payload_addr,
      io_input_arw_payload_len => dbus_axi_arw_payload_len,
      io_input_arw_payload_size => dbus_axi_arw_payload_size,
      io_input_arw_payload_cache => dbus_axi_arw_payload_cache,
      io_input_arw_payload_prot => dbus_axi_arw_payload_prot,
      io_input_arw_payload_write => dbus_axi_arw_payload_write,
      io_input_w_valid => dbus_axi_w_valid,
      io_input_w_ready => dbus_axi_decoder_io_input_w_ready,
      io_input_w_payload_data => dbus_axi_w_payload_data,
      io_input_w_payload_strb => dbus_axi_w_payload_strb,
      io_input_w_payload_last => dbus_axi_w_payload_last,
      io_input_b_valid => dbus_axi_decoder_io_input_b_valid,
      io_input_b_ready => dbus_axi_b_ready,
      io_input_b_payload_resp => dbus_axi_decoder_io_input_b_payload_resp,
      io_input_r_valid => dbus_axi_decoder_io_input_r_valid,
      io_input_r_ready => dbus_axi_decoder_io_input_r_ready,
      io_input_r_payload_data => dbus_axi_decoder_io_input_r_payload_data,
      io_input_r_payload_resp => dbus_axi_decoder_io_input_r_payload_resp,
      io_input_r_payload_last => dbus_axi_decoder_io_input_r_payload_last,
      io_sharedOutputs_0_arw_valid => dbus_axi_decoder_io_sharedOutputs_0_arw_valid,
      io_sharedOutputs_0_arw_ready => dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_fire_1,
      io_sharedOutputs_0_arw_payload_addr => dbus_axi_decoder_io_sharedOutputs_0_arw_payload_addr,
      io_sharedOutputs_0_arw_payload_len => dbus_axi_decoder_io_sharedOutputs_0_arw_payload_len,
      io_sharedOutputs_0_arw_payload_size => dbus_axi_decoder_io_sharedOutputs_0_arw_payload_size,
      io_sharedOutputs_0_arw_payload_cache => dbus_axi_decoder_io_sharedOutputs_0_arw_payload_cache,
      io_sharedOutputs_0_arw_payload_prot => dbus_axi_decoder_io_sharedOutputs_0_arw_payload_prot,
      io_sharedOutputs_0_arw_payload_write => dbus_axi_decoder_io_sharedOutputs_0_arw_payload_write,
      io_sharedOutputs_0_w_valid => dbus_axi_decoder_io_sharedOutputs_0_w_valid,
      io_sharedOutputs_0_w_ready => axi_ram_io_axi_arbiter_io_sharedInputs_0_w_ready,
      io_sharedOutputs_0_w_payload_data => dbus_axi_decoder_io_sharedOutputs_0_w_payload_data,
      io_sharedOutputs_0_w_payload_strb => dbus_axi_decoder_io_sharedOutputs_0_w_payload_strb,
      io_sharedOutputs_0_w_payload_last => dbus_axi_decoder_io_sharedOutputs_0_w_payload_last,
      io_sharedOutputs_0_b_valid => axi_ram_io_axi_arbiter_io_sharedInputs_0_b_valid,
      io_sharedOutputs_0_b_ready => dbus_axi_decoder_io_sharedOutputs_0_b_ready,
      io_sharedOutputs_0_b_payload_resp => axi_ram_io_axi_arbiter_io_sharedInputs_0_b_payload_resp,
      io_sharedOutputs_0_r_valid => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_valid,
      io_sharedOutputs_0_r_ready => dbus_axi_decoder_io_sharedOutputs_0_r_ready,
      io_sharedOutputs_0_r_payload_data => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_data,
      io_sharedOutputs_0_r_payload_resp => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_resp,
      io_sharedOutputs_0_r_payload_last => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_last,
      io_sharedOutputs_1_arw_valid => dbus_axi_decoder_io_sharedOutputs_1_arw_valid,
      io_sharedOutputs_1_arw_ready => dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_fire_1,
      io_sharedOutputs_1_arw_payload_addr => dbus_axi_decoder_io_sharedOutputs_1_arw_payload_addr,
      io_sharedOutputs_1_arw_payload_len => dbus_axi_decoder_io_sharedOutputs_1_arw_payload_len,
      io_sharedOutputs_1_arw_payload_size => dbus_axi_decoder_io_sharedOutputs_1_arw_payload_size,
      io_sharedOutputs_1_arw_payload_cache => dbus_axi_decoder_io_sharedOutputs_1_arw_payload_cache,
      io_sharedOutputs_1_arw_payload_prot => dbus_axi_decoder_io_sharedOutputs_1_arw_payload_prot,
      io_sharedOutputs_1_arw_payload_write => dbus_axi_decoder_io_sharedOutputs_1_arw_payload_write,
      io_sharedOutputs_1_w_valid => dbus_axi_decoder_io_sharedOutputs_1_w_valid,
      io_sharedOutputs_1_w_ready => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_w_ready,
      io_sharedOutputs_1_w_payload_data => dbus_axi_decoder_io_sharedOutputs_1_w_payload_data,
      io_sharedOutputs_1_w_payload_strb => dbus_axi_decoder_io_sharedOutputs_1_w_payload_strb,
      io_sharedOutputs_1_w_payload_last => dbus_axi_decoder_io_sharedOutputs_1_w_payload_last,
      io_sharedOutputs_1_b_valid => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_valid,
      io_sharedOutputs_1_b_ready => dbus_axi_decoder_io_sharedOutputs_1_b_ready,
      io_sharedOutputs_1_b_payload_resp => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_payload_resp,
      io_sharedOutputs_1_r_valid => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_valid,
      io_sharedOutputs_1_r_ready => dbus_axi_decoder_io_sharedOutputs_1_r_ready,
      io_sharedOutputs_1_r_payload_data => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_data,
      io_sharedOutputs_1_r_payload_resp => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_resp,
      io_sharedOutputs_1_r_payload_last => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_ram_io_axi_arbiter : entity work.Axi4SharedArbiter
    port map ( 
      io_readInputs_0_ar_valid => axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_valid,
      io_readInputs_0_ar_ready => axi_ram_io_axi_arbiter_io_readInputs_0_ar_ready,
      io_readInputs_0_ar_payload_addr => axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr,
      io_readInputs_0_ar_payload_id => zz_io_readInputs_0_ar_payload_id,
      io_readInputs_0_ar_payload_len => axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_len,
      io_readInputs_0_ar_payload_size => pkg_unsigned("010"),
      io_readInputs_0_ar_payload_burst => axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_burst,
      io_readInputs_0_r_valid => axi_ram_io_axi_arbiter_io_readInputs_0_r_valid,
      io_readInputs_0_r_ready => axi4ReadOnlyDecoder_1_io_outputs_0_r_ready,
      io_readInputs_0_r_payload_data => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_data,
      io_readInputs_0_r_payload_id => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_id,
      io_readInputs_0_r_payload_resp => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_resp,
      io_readInputs_0_r_payload_last => axi_ram_io_axi_arbiter_io_readInputs_0_r_payload_last,
      io_sharedInputs_0_arw_valid => dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_valid,
      io_sharedInputs_0_arw_ready => axi_ram_io_axi_arbiter_io_sharedInputs_0_arw_ready,
      io_sharedInputs_0_arw_payload_addr => axi_ram_io_axi_arbiter_io_sharedInputs_0_arw_payload_addr,
      io_sharedInputs_0_arw_payload_id => zz_io_sharedInputs_0_arw_payload_id,
      io_sharedInputs_0_arw_payload_len => dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_len,
      io_sharedInputs_0_arw_payload_size => dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_size,
      io_sharedInputs_0_arw_payload_burst => pkg_stdLogicVector("01"),
      io_sharedInputs_0_arw_payload_write => dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_write,
      io_sharedInputs_0_w_valid => dbus_axi_decoder_io_sharedOutputs_0_w_valid,
      io_sharedInputs_0_w_ready => axi_ram_io_axi_arbiter_io_sharedInputs_0_w_ready,
      io_sharedInputs_0_w_payload_data => dbus_axi_decoder_io_sharedOutputs_0_w_payload_data,
      io_sharedInputs_0_w_payload_strb => dbus_axi_decoder_io_sharedOutputs_0_w_payload_strb,
      io_sharedInputs_0_w_payload_last => dbus_axi_decoder_io_sharedOutputs_0_w_payload_last,
      io_sharedInputs_0_b_valid => axi_ram_io_axi_arbiter_io_sharedInputs_0_b_valid,
      io_sharedInputs_0_b_ready => dbus_axi_decoder_io_sharedOutputs_0_b_ready,
      io_sharedInputs_0_b_payload_id => axi_ram_io_axi_arbiter_io_sharedInputs_0_b_payload_id,
      io_sharedInputs_0_b_payload_resp => axi_ram_io_axi_arbiter_io_sharedInputs_0_b_payload_resp,
      io_sharedInputs_0_r_valid => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_valid,
      io_sharedInputs_0_r_ready => dbus_axi_decoder_io_sharedOutputs_0_r_ready,
      io_sharedInputs_0_r_payload_data => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_data,
      io_sharedInputs_0_r_payload_id => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_id,
      io_sharedInputs_0_r_payload_resp => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_resp,
      io_sharedInputs_0_r_payload_last => axi_ram_io_axi_arbiter_io_sharedInputs_0_r_payload_last,
      io_output_arw_valid => axi_ram_io_axi_arbiter_io_output_arw_valid,
      io_output_arw_ready => axi_ram_io_axi_arbiter_io_output_arw_ready,
      io_output_arw_payload_addr => axi_ram_io_axi_arbiter_io_output_arw_payload_addr,
      io_output_arw_payload_id => axi_ram_io_axi_arbiter_io_output_arw_payload_id,
      io_output_arw_payload_len => axi_ram_io_axi_arbiter_io_output_arw_payload_len,
      io_output_arw_payload_size => axi_ram_io_axi_arbiter_io_output_arw_payload_size,
      io_output_arw_payload_burst => axi_ram_io_axi_arbiter_io_output_arw_payload_burst,
      io_output_arw_payload_write => axi_ram_io_axi_arbiter_io_output_arw_payload_write,
      io_output_w_valid => axi_ram_io_axi_arbiter_io_output_w_valid,
      io_output_w_ready => axi_ram_io_axi_arbiter_io_output_w_ready,
      io_output_w_payload_data => axi_ram_io_axi_arbiter_io_output_w_payload_data,
      io_output_w_payload_strb => axi_ram_io_axi_arbiter_io_output_w_payload_strb,
      io_output_w_payload_last => axi_ram_io_axi_arbiter_io_output_w_payload_last,
      io_output_b_valid => axi_ram_io_axi_b_valid,
      io_output_b_ready => axi_ram_io_axi_arbiter_io_output_b_ready,
      io_output_b_payload_id => axi_ram_io_axi_b_payload_id,
      io_output_b_payload_resp => axi_ram_io_axi_b_payload_resp,
      io_output_r_valid => axi_ram_io_axi_r_valid,
      io_output_r_ready => axi_ram_io_axi_arbiter_io_output_r_ready,
      io_output_r_payload_data => axi_ram_io_axi_r_payload_data,
      io_output_r_payload_id => axi_ram_io_axi_r_payload_id,
      io_output_r_payload_resp => axi_ram_io_axi_r_payload_resp,
      io_output_r_payload_last => axi_ram_io_axi_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  axi_apbBridge_io_axi_arbiter : entity work.Axi4SharedArbiter_1
    port map ( 
      io_sharedInputs_0_arw_valid => dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_valid,
      io_sharedInputs_0_arw_ready => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_arw_ready,
      io_sharedInputs_0_arw_payload_addr => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_arw_payload_addr,
      io_sharedInputs_0_arw_payload_id => zz_io_sharedInputs_0_arw_payload_id_1,
      io_sharedInputs_0_arw_payload_len => dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_len,
      io_sharedInputs_0_arw_payload_size => dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_size,
      io_sharedInputs_0_arw_payload_burst => pkg_stdLogicVector("01"),
      io_sharedInputs_0_arw_payload_write => dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_write,
      io_sharedInputs_0_w_valid => dbus_axi_decoder_io_sharedOutputs_1_w_valid,
      io_sharedInputs_0_w_ready => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_w_ready,
      io_sharedInputs_0_w_payload_data => dbus_axi_decoder_io_sharedOutputs_1_w_payload_data,
      io_sharedInputs_0_w_payload_strb => dbus_axi_decoder_io_sharedOutputs_1_w_payload_strb,
      io_sharedInputs_0_w_payload_last => dbus_axi_decoder_io_sharedOutputs_1_w_payload_last,
      io_sharedInputs_0_b_valid => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_valid,
      io_sharedInputs_0_b_ready => dbus_axi_decoder_io_sharedOutputs_1_b_ready,
      io_sharedInputs_0_b_payload_id => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_payload_id,
      io_sharedInputs_0_b_payload_resp => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_b_payload_resp,
      io_sharedInputs_0_r_valid => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_valid,
      io_sharedInputs_0_r_ready => dbus_axi_decoder_io_sharedOutputs_1_r_ready,
      io_sharedInputs_0_r_payload_data => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_data,
      io_sharedInputs_0_r_payload_id => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_id,
      io_sharedInputs_0_r_payload_resp => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_resp,
      io_sharedInputs_0_r_payload_last => axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_r_payload_last,
      io_output_arw_valid => axi_apbBridge_io_axi_arbiter_io_output_arw_valid,
      io_output_arw_ready => axi_apbBridge_io_axi_arbiter_io_output_arw_ready,
      io_output_arw_payload_addr => axi_apbBridge_io_axi_arbiter_io_output_arw_payload_addr,
      io_output_arw_payload_id => axi_apbBridge_io_axi_arbiter_io_output_arw_payload_id,
      io_output_arw_payload_len => axi_apbBridge_io_axi_arbiter_io_output_arw_payload_len,
      io_output_arw_payload_size => axi_apbBridge_io_axi_arbiter_io_output_arw_payload_size,
      io_output_arw_payload_burst => axi_apbBridge_io_axi_arbiter_io_output_arw_payload_burst,
      io_output_arw_payload_write => axi_apbBridge_io_axi_arbiter_io_output_arw_payload_write,
      io_output_w_valid => axi_apbBridge_io_axi_arbiter_io_output_w_valid,
      io_output_w_ready => axi_apbBridge_io_axi_arbiter_io_output_w_ready,
      io_output_w_payload_data => axi_apbBridge_io_axi_arbiter_io_output_w_payload_data,
      io_output_w_payload_strb => axi_apbBridge_io_axi_arbiter_io_output_w_payload_strb,
      io_output_w_payload_last => axi_apbBridge_io_axi_arbiter_io_output_w_payload_last,
      io_output_b_valid => axi_apbBridge_io_axi_b_valid,
      io_output_b_ready => axi_apbBridge_io_axi_arbiter_io_output_b_ready,
      io_output_b_payload_id => axi_apbBridge_io_axi_b_payload_id,
      io_output_b_payload_resp => axi_apbBridge_io_axi_b_payload_resp,
      io_output_r_valid => axi_apbBridge_io_axi_r_valid,
      io_output_r_ready => axi_apbBridge_io_axi_arbiter_io_output_r_ready,
      io_output_r_payload_data => axi_apbBridge_io_axi_r_payload_data,
      io_output_r_payload_id => axi_apbBridge_io_axi_r_payload_id,
      io_output_r_payload_resp => axi_apbBridge_io_axi_r_payload_resp,
      io_output_r_payload_last => axi_apbBridge_io_axi_r_payload_last,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  io_apb_decoder : entity work.Apb3Decoder
    port map ( 
      io_input_PADDR => axi_apbBridge_io_apb_PADDR,
      io_input_PSEL => axi_apbBridge_io_apb_PSEL,
      io_input_PENABLE => axi_apbBridge_io_apb_PENABLE,
      io_input_PREADY => io_apb_decoder_io_input_PREADY,
      io_input_PWRITE => axi_apbBridge_io_apb_PWRITE,
      io_input_PWDATA => axi_apbBridge_io_apb_PWDATA,
      io_input_PRDATA => io_apb_decoder_io_input_PRDATA,
      io_input_PSLVERROR => io_apb_decoder_io_input_PSLVERROR,
      io_output_PADDR => io_apb_decoder_io_output_PADDR,
      io_output_PSEL => io_apb_decoder_io_output_PSEL,
      io_output_PENABLE => io_apb_decoder_io_output_PENABLE,
      io_output_PREADY => apb3Router_1_io_input_PREADY,
      io_output_PWRITE => io_apb_decoder_io_output_PWRITE,
      io_output_PWDATA => io_apb_decoder_io_output_PWDATA,
      io_output_PRDATA => apb3Router_1_io_input_PRDATA,
      io_output_PSLVERROR => apb3Router_1_io_input_PSLVERROR 
    );
  apb3Router_1 : entity work.Apb3Router
    port map ( 
      io_input_PADDR => io_apb_decoder_io_output_PADDR,
      io_input_PSEL => io_apb_decoder_io_output_PSEL,
      io_input_PENABLE => io_apb_decoder_io_output_PENABLE,
      io_input_PREADY => apb3Router_1_io_input_PREADY,
      io_input_PWRITE => io_apb_decoder_io_output_PWRITE,
      io_input_PWDATA => io_apb_decoder_io_output_PWDATA,
      io_input_PRDATA => apb3Router_1_io_input_PRDATA,
      io_input_PSLVERROR => apb3Router_1_io_input_PSLVERROR,
      io_outputs_0_PADDR => apb3Router_1_io_outputs_0_PADDR,
      io_outputs_0_PSEL => apb3Router_1_io_outputs_0_PSEL,
      io_outputs_0_PENABLE => apb3Router_1_io_outputs_0_PENABLE,
      io_outputs_0_PREADY => axi_gpioACtrl_io_apb_PREADY,
      io_outputs_0_PWRITE => apb3Router_1_io_outputs_0_PWRITE,
      io_outputs_0_PWDATA => apb3Router_1_io_outputs_0_PWDATA,
      io_outputs_0_PRDATA => axi_gpioACtrl_io_apb_PRDATA,
      io_outputs_0_PSLVERROR => axi_gpioACtrl_io_apb_PSLVERROR,
      io_outputs_1_PADDR => apb3Router_1_io_outputs_1_PADDR,
      io_outputs_1_PSEL => apb3Router_1_io_outputs_1_PSEL,
      io_outputs_1_PENABLE => apb3Router_1_io_outputs_1_PENABLE,
      io_outputs_1_PREADY => axi_uartCtrl_io_apb_PREADY,
      io_outputs_1_PWRITE => apb3Router_1_io_outputs_1_PWRITE,
      io_outputs_1_PWDATA => apb3Router_1_io_outputs_1_PWDATA,
      io_outputs_1_PRDATA => axi_uartCtrl_io_apb_PRDATA,
      io_outputs_1_PSLVERROR => pkg_toStdLogic(false),
      io_outputs_2_PADDR => apb3Router_1_io_outputs_2_PADDR,
      io_outputs_2_PSEL => apb3Router_1_io_outputs_2_PSEL,
      io_outputs_2_PENABLE => apb3Router_1_io_outputs_2_PENABLE,
      io_outputs_2_PREADY => axi_timer_io_apb_PREADY,
      io_outputs_2_PWRITE => apb3Router_1_io_outputs_2_PWRITE,
      io_outputs_2_PWDATA => apb3Router_1_io_outputs_2_PWDATA,
      io_outputs_2_PRDATA => axi_timer_io_apb_PRDATA,
      io_outputs_2_PSLVERROR => axi_timer_io_apb_PSLVERROR,
      io_mainClk => io_mainClk,
      resetCtrl_axiReset => resetCtrl_axiReset 
    );
  process(when_Muraxy_l198)
  begin
    resetCtrl_systemResetUnbuffered <= pkg_toStdLogic(false);
    if when_Muraxy_l198 = '1' then
      resetCtrl_systemResetUnbuffered <= pkg_toStdLogic(true);
    end if;
  end process;

  zz_when_Muraxy_l198(5 downto 0) <= pkg_unsigned("111111");
  when_Muraxy_l198 <= pkg_toStdLogic(resetCtrl_systemResetCounter /= zz_when_Muraxy_l198);
  when_Muraxy_l202 <= io_asyncReset_buffercc_io_dataOut;
  axi_core_cpu_iBus_rsp_payload_error <= (not pkg_toStdLogic(axi4ReadOnlyDecoder_1_io_input_r_payload_resp = pkg_stdLogicVector("00")));
  process(axi_core_cpu_dBus_cmd_m2sPipe_ready,when_Stream_l342)
  begin
    axi_core_cpu_dBus_cmd_ready <= axi_core_cpu_dBus_cmd_m2sPipe_ready;
    if when_Stream_l342 = '1' then
      axi_core_cpu_dBus_cmd_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Stream_l342 <= (not axi_core_cpu_dBus_cmd_m2sPipe_valid);
  axi_core_cpu_dBus_cmd_m2sPipe_valid <= axi_core_cpu_dBus_cmd_rValid;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_wr <= axi_core_cpu_dBus_cmd_rData_wr;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_uncached <= axi_core_cpu_dBus_cmd_rData_uncached;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_address <= axi_core_cpu_dBus_cmd_rData_address;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_data <= axi_core_cpu_dBus_cmd_rData_data;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_mask <= axi_core_cpu_dBus_cmd_rData_mask;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_size <= axi_core_cpu_dBus_cmd_rData_size;
  axi_core_cpu_dBus_cmd_m2sPipe_payload_last <= axi_core_cpu_dBus_cmd_rData_last;
  process(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_ready,when_Stream_l342_1)
  begin
    axi_core_cpu_dBus_cmd_m2sPipe_ready <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_ready;
    if when_Stream_l342_1 = '1' then
      axi_core_cpu_dBus_cmd_m2sPipe_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Stream_l342_1 <= (not axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_valid);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_valid <= axi_core_cpu_dBus_cmd_m2sPipe_rValid;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_wr <= axi_core_cpu_dBus_cmd_m2sPipe_rData_wr;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_uncached <= axi_core_cpu_dBus_cmd_m2sPipe_rData_uncached;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_address <= axi_core_cpu_dBus_cmd_m2sPipe_rData_address;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_data <= axi_core_cpu_dBus_cmd_m2sPipe_rData_data;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_mask <= axi_core_cpu_dBus_cmd_m2sPipe_rData_mask;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_size <= axi_core_cpu_dBus_cmd_m2sPipe_rData_size;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_last <= axi_core_cpu_dBus_cmd_m2sPipe_rData_last;
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_ready <= (not axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_valid <= (axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_valid or axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_wr <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_wr,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_wr);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_uncached <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_uncached,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_uncached);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_address <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_address,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_address);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_data <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_data,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_data);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_mask <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_mask,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_mask);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_size <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_size,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_size);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_last <= pkg_mux(axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_last,axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_last);
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_fire <= (axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_valid and axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready);
  when_Utils_l594 <= (axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_fire and axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_wr);
  dbus_axi_b_fire <= (dbus_axi_b_valid and dbus_axi_b_ready);
  process(when_Utils_l594)
  begin
    zz_when_Utils_l622 <= pkg_toStdLogic(false);
    if when_Utils_l594 = '1' then
      zz_when_Utils_l622 <= pkg_toStdLogic(true);
    end if;
  end process;

  process(dbus_axi_b_fire)
  begin
    zz_when_Utils_l622_1 <= pkg_toStdLogic(false);
    if dbus_axi_b_fire = '1' then
      zz_when_Utils_l622_1 <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Utils_l622 <= (zz_when_Utils_l622 and (not zz_when_Utils_l622_1));
  process(when_Utils_l622,when_Utils_l624)
  begin
    if when_Utils_l622 = '1' then
      zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_1 <= pkg_unsigned("001");
    else
      if when_Utils_l624 = '1' then
        zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_1 <= pkg_unsigned("111");
      else
        zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_1 <= pkg_unsigned("000");
      end if;
    end if;
  end process;

  when_Utils_l624 <= ((not zz_when_Utils_l622) and zz_when_Utils_l622_1);
  zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_2 <= (not ((pkg_toStdLogic(zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready /= pkg_unsigned("000")) and (not axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_payload_wr)) or pkg_toStdLogic(zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready = pkg_unsigned("111"))));
  axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready <= (streamFork_3_io_input_ready and zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_2);
  streamFork_3_io_input_valid <= (axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_valid and zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_2);
  streamFork_3_io_outputs_0_fire <= (streamFork_3_io_outputs_0_valid and streamFork_3_io_outputs_0_ready);
  process(streamFork_3_io_outputs_0_valid,zz_1)
  begin
    streamFork_3_io_outputs_0_thrown_valid <= streamFork_3_io_outputs_0_valid;
    if zz_1 = '1' then
      streamFork_3_io_outputs_0_thrown_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  process(streamFork_3_io_outputs_0_thrown_ready,zz_1)
  begin
    streamFork_3_io_outputs_0_ready <= streamFork_3_io_outputs_0_thrown_ready;
    if zz_1 = '1' then
      streamFork_3_io_outputs_0_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  streamFork_3_io_outputs_0_thrown_payload_wr <= streamFork_3_io_outputs_0_payload_wr;
  streamFork_3_io_outputs_0_thrown_payload_uncached <= streamFork_3_io_outputs_0_payload_uncached;
  streamFork_3_io_outputs_0_thrown_payload_address <= streamFork_3_io_outputs_0_payload_address;
  streamFork_3_io_outputs_0_thrown_payload_data <= streamFork_3_io_outputs_0_payload_data;
  streamFork_3_io_outputs_0_thrown_payload_mask <= streamFork_3_io_outputs_0_payload_mask;
  streamFork_3_io_outputs_0_thrown_payload_size <= streamFork_3_io_outputs_0_payload_size;
  streamFork_3_io_outputs_0_thrown_payload_last <= streamFork_3_io_outputs_0_payload_last;
  when_Stream_l408 <= (not streamFork_3_io_outputs_1_payload_wr);
  process(streamFork_3_io_outputs_1_valid,when_Stream_l408)
  begin
    streamFork_3_io_outputs_1_thrown_valid <= streamFork_3_io_outputs_1_valid;
    if when_Stream_l408 = '1' then
      streamFork_3_io_outputs_1_thrown_valid <= pkg_toStdLogic(false);
    end if;
  end process;

  process(streamFork_3_io_outputs_1_thrown_ready,when_Stream_l408)
  begin
    streamFork_3_io_outputs_1_ready <= streamFork_3_io_outputs_1_thrown_ready;
    if when_Stream_l408 = '1' then
      streamFork_3_io_outputs_1_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  streamFork_3_io_outputs_1_thrown_payload_wr <= streamFork_3_io_outputs_1_payload_wr;
  streamFork_3_io_outputs_1_thrown_payload_uncached <= streamFork_3_io_outputs_1_payload_uncached;
  streamFork_3_io_outputs_1_thrown_payload_address <= streamFork_3_io_outputs_1_payload_address;
  streamFork_3_io_outputs_1_thrown_payload_data <= streamFork_3_io_outputs_1_payload_data;
  streamFork_3_io_outputs_1_thrown_payload_mask <= streamFork_3_io_outputs_1_payload_mask;
  streamFork_3_io_outputs_1_thrown_payload_size <= streamFork_3_io_outputs_1_payload_size;
  streamFork_3_io_outputs_1_thrown_payload_last <= streamFork_3_io_outputs_1_payload_last;
  dbus_axi_arw_valid <= streamFork_3_io_outputs_0_thrown_valid;
  streamFork_3_io_outputs_0_thrown_ready <= dbus_axi_arw_ready;
  dbus_axi_arw_payload_write <= streamFork_3_io_outputs_0_thrown_payload_wr;
  dbus_axi_arw_payload_prot <= pkg_stdLogicVector("010");
  dbus_axi_arw_payload_cache <= pkg_stdLogicVector("1111");
  dbus_axi_arw_payload_size <= pkg_unsigned("010");
  dbus_axi_arw_payload_addr <= streamFork_3_io_outputs_0_thrown_payload_address;
  dbus_axi_arw_payload_len <= pkg_resize(pkg_mux(pkg_toStdLogic(streamFork_3_io_outputs_0_thrown_payload_size = pkg_unsigned("101")),pkg_unsigned("111"),pkg_unsigned("000")),8);
  dbus_axi_w_valid <= streamFork_3_io_outputs_1_thrown_valid;
  streamFork_3_io_outputs_1_thrown_ready <= dbus_axi_w_ready;
  dbus_axi_w_payload_data <= streamFork_3_io_outputs_1_thrown_payload_data;
  dbus_axi_w_payload_strb <= streamFork_3_io_outputs_1_thrown_payload_mask;
  dbus_axi_w_payload_last <= streamFork_3_io_outputs_1_thrown_payload_last;
  axi_core_cpu_dBus_rsp_payload_error <= (not pkg_toStdLogic(dbus_axi_r_payload_resp = pkg_stdLogicVector("00")));
  dbus_axi_r_ready <= pkg_toStdLogic(true);
  dbus_axi_b_ready <= pkg_toStdLogic(true);
  axi_core_cpu_debug_bus_cmd_payload_address <= pkg_resize(systemDebugger_1_io_mem_cmd_payload_address,8);
  axi_core_cpu_debug_bus_cmd_fire <= (systemDebugger_1_io_mem_cmd_valid and axi_core_cpu_debug_bus_cmd_ready);
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_fire <= (axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_valid and axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_ready);
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_fire_1 <= (axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_valid and axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_ready);
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_valid <= axi4ReadOnlyDecoder_1_io_outputs_0_ar_rValid;
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_addr <= axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_addr;
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_len <= axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_len;
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_burst <= axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_burst;
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_cache <= axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_cache;
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_prot <= axi4ReadOnlyDecoder_1_io_outputs_0_ar_payload_prot;
  axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_ready <= axi_ram_io_axi_arbiter_io_readInputs_0_ar_ready;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_fire <= (dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_valid and dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_ready);
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_fire_1 <= (dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_valid and dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_ready);
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_valid <= dbus_axi_decoder_io_sharedOutputs_0_arw_rValid;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_addr <= dbus_axi_decoder_io_sharedOutputs_0_arw_payload_addr;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_len <= dbus_axi_decoder_io_sharedOutputs_0_arw_payload_len;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_size <= dbus_axi_decoder_io_sharedOutputs_0_arw_payload_size;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_cache <= dbus_axi_decoder_io_sharedOutputs_0_arw_payload_cache;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_prot <= dbus_axi_decoder_io_sharedOutputs_0_arw_payload_prot;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_write <= dbus_axi_decoder_io_sharedOutputs_0_arw_payload_write;
  dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_ready <= axi_ram_io_axi_arbiter_io_sharedInputs_0_arw_ready;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_fire <= (dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_valid and dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_ready);
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_fire_1 <= (dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_valid and dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_ready);
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_valid <= dbus_axi_decoder_io_sharedOutputs_1_arw_rValid;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_addr <= dbus_axi_decoder_io_sharedOutputs_1_arw_payload_addr;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_len <= dbus_axi_decoder_io_sharedOutputs_1_arw_payload_len;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_size <= dbus_axi_decoder_io_sharedOutputs_1_arw_payload_size;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_cache <= dbus_axi_decoder_io_sharedOutputs_1_arw_payload_cache;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_prot <= dbus_axi_decoder_io_sharedOutputs_1_arw_payload_prot;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_write <= dbus_axi_decoder_io_sharedOutputs_1_arw_payload_write;
  dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_ready <= axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_arw_ready;
  dbus_axi_arw_ready <= dbus_axi_decoder_io_input_arw_ready;
  dbus_axi_w_ready <= dbus_axi_decoder_io_input_w_ready;
  dbus_axi_b_valid <= dbus_axi_decoder_io_input_b_valid;
  dbus_axi_b_payload_resp <= dbus_axi_decoder_io_input_b_payload_resp;
  process(dbus_axi_decoder_io_input_r_m2sPipe_ready,when_Stream_l342_2)
  begin
    dbus_axi_decoder_io_input_r_ready <= dbus_axi_decoder_io_input_r_m2sPipe_ready;
    if when_Stream_l342_2 = '1' then
      dbus_axi_decoder_io_input_r_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Stream_l342_2 <= (not dbus_axi_decoder_io_input_r_m2sPipe_valid);
  dbus_axi_decoder_io_input_r_m2sPipe_valid <= dbus_axi_decoder_io_input_r_rValid;
  dbus_axi_decoder_io_input_r_m2sPipe_payload_data <= dbus_axi_decoder_io_input_r_rData_data;
  dbus_axi_decoder_io_input_r_m2sPipe_payload_resp <= dbus_axi_decoder_io_input_r_rData_resp;
  dbus_axi_decoder_io_input_r_m2sPipe_payload_last <= dbus_axi_decoder_io_input_r_rData_last;
  dbus_axi_r_valid <= dbus_axi_decoder_io_input_r_m2sPipe_valid;
  dbus_axi_decoder_io_input_r_m2sPipe_ready <= dbus_axi_r_ready;
  dbus_axi_r_payload_data <= dbus_axi_decoder_io_input_r_m2sPipe_payload_data;
  dbus_axi_r_payload_resp <= dbus_axi_decoder_io_input_r_m2sPipe_payload_resp;
  dbus_axi_r_payload_last <= dbus_axi_decoder_io_input_r_m2sPipe_payload_last;
  axi_ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr <= pkg_resize(axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_payload_addr,15);
  zz_io_readInputs_0_ar_payload_id(2 downto 0) <= pkg_unsigned("000");
  axi_ram_io_axi_arbiter_io_sharedInputs_0_arw_payload_addr <= pkg_resize(dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_payload_addr,15);
  zz_io_sharedInputs_0_arw_payload_id(2 downto 0) <= pkg_unsigned("000");
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_fire <= (axi_ram_io_axi_arbiter_io_output_arw_halfPipe_valid and axi_ram_io_axi_arbiter_io_output_arw_halfPipe_ready);
  axi_ram_io_axi_arbiter_io_output_arw_ready <= (not axi_ram_io_axi_arbiter_io_output_arw_rValid);
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_valid <= axi_ram_io_axi_arbiter_io_output_arw_rValid;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_addr <= axi_ram_io_axi_arbiter_io_output_arw_rData_addr;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_id <= axi_ram_io_axi_arbiter_io_output_arw_rData_id;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_len <= axi_ram_io_axi_arbiter_io_output_arw_rData_len;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_size <= axi_ram_io_axi_arbiter_io_output_arw_rData_size;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_burst <= axi_ram_io_axi_arbiter_io_output_arw_rData_burst;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_payload_write <= axi_ram_io_axi_arbiter_io_output_arw_rData_write;
  axi_ram_io_axi_arbiter_io_output_arw_halfPipe_ready <= axi_ram_io_axi_arw_ready;
  axi_ram_io_axi_arbiter_io_output_w_ready <= (not axi_ram_io_axi_arbiter_io_output_w_rValid);
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_valid <= (axi_ram_io_axi_arbiter_io_output_w_valid or axi_ram_io_axi_arbiter_io_output_w_rValid);
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_data <= pkg_mux(axi_ram_io_axi_arbiter_io_output_w_rValid,axi_ram_io_axi_arbiter_io_output_w_rData_data,axi_ram_io_axi_arbiter_io_output_w_payload_data);
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_strb <= pkg_mux(axi_ram_io_axi_arbiter_io_output_w_rValid,axi_ram_io_axi_arbiter_io_output_w_rData_strb,axi_ram_io_axi_arbiter_io_output_w_payload_strb);
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_last <= pkg_mux(axi_ram_io_axi_arbiter_io_output_w_rValid,axi_ram_io_axi_arbiter_io_output_w_rData_last,axi_ram_io_axi_arbiter_io_output_w_payload_last);
  process(axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_ready,when_Stream_l342_3)
  begin
    axi_ram_io_axi_arbiter_io_output_w_s2mPipe_ready <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_ready;
    if when_Stream_l342_3 = '1' then
      axi_ram_io_axi_arbiter_io_output_w_s2mPipe_ready <= pkg_toStdLogic(true);
    end if;
  end process;

  when_Stream_l342_3 <= (not axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_valid);
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_valid <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rValid;
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_data <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_data;
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_strb <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_strb;
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_payload_last <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_last;
  axi_ram_io_axi_arbiter_io_output_w_s2mPipe_m2sPipe_ready <= axi_ram_io_axi_w_ready;
  axi_apbBridge_io_axi_arbiter_io_sharedInputs_0_arw_payload_addr <= pkg_resize(dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_payload_addr,20);
  zz_io_sharedInputs_0_arw_payload_id_1(3 downto 0) <= pkg_unsigned("0000");
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_fire <= (axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_valid and axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_ready);
  axi_apbBridge_io_axi_arbiter_io_output_arw_ready <= (not axi_apbBridge_io_axi_arbiter_io_output_arw_rValid);
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_valid <= axi_apbBridge_io_axi_arbiter_io_output_arw_rValid;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_addr <= axi_apbBridge_io_axi_arbiter_io_output_arw_rData_addr;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_id <= axi_apbBridge_io_axi_arbiter_io_output_arw_rData_id;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_len <= axi_apbBridge_io_axi_arbiter_io_output_arw_rData_len;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_size <= axi_apbBridge_io_axi_arbiter_io_output_arw_rData_size;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_burst <= axi_apbBridge_io_axi_arbiter_io_output_arw_rData_burst;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_payload_write <= axi_apbBridge_io_axi_arbiter_io_output_arw_rData_write;
  axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_ready <= axi_apbBridge_io_axi_arw_ready;
  axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_fire <= (axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_valid and axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_ready);
  axi_apbBridge_io_axi_arbiter_io_output_w_ready <= (not axi_apbBridge_io_axi_arbiter_io_output_w_rValid);
  axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_valid <= axi_apbBridge_io_axi_arbiter_io_output_w_rValid;
  axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_data <= axi_apbBridge_io_axi_arbiter_io_output_w_rData_data;
  axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_strb <= axi_apbBridge_io_axi_arbiter_io_output_w_rData_strb;
  axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_payload_last <= axi_apbBridge_io_axi_arbiter_io_output_w_rData_last;
  axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_ready <= axi_apbBridge_io_axi_w_ready;
  axi_gpioACtrl_io_apb_PADDR <= pkg_resize(apb3Router_1_io_outputs_0_PADDR,4);
  axi_uartCtrl_io_apb_PADDR <= pkg_resize(apb3Router_1_io_outputs_1_PADDR,5);
  axi_timer_io_apb_PADDR <= pkg_resize(apb3Router_1_io_outputs_2_PADDR,8);
  io_gpioA_write <= axi_gpioACtrl_io_gpio_write;
  io_gpioA_writeEnable <= axi_gpioACtrl_io_gpio_writeEnable;
  io_uart_txd <= axi_uartCtrl_io_uart_txd;
  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if when_Muraxy_l198 = '1' then
        resetCtrl_systemResetCounter <= (resetCtrl_systemResetCounter + pkg_unsigned("000001"));
      end if;
      if when_Muraxy_l202 = '1' then
        resetCtrl_systemResetCounter <= pkg_unsigned("000000");
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      resetCtrl_systemReset <= resetCtrl_systemResetUnbuffered;
      resetCtrl_axiReset <= resetCtrl_systemResetUnbuffered;
      if axi_core_cpu_debug_resetOut_regNext = '1' then
        resetCtrl_axiReset <= pkg_toStdLogic(true);
      end if;
    end if;
  end process;

  process(io_mainClk, resetCtrl_axiReset)
  begin
    if resetCtrl_axiReset = '1' then
      axi_core_cpu_dBus_cmd_rValid <= pkg_toStdLogic(false);
      axi_core_cpu_dBus_cmd_m2sPipe_rValid <= pkg_toStdLogic(false);
      axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid <= pkg_toStdLogic(false);
      zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready <= pkg_unsigned("000");
      zz_1 <= pkg_toStdLogic(false);
      axi4ReadOnlyDecoder_1_io_outputs_0_ar_rValid <= pkg_toStdLogic(false);
      dbus_axi_decoder_io_sharedOutputs_0_arw_rValid <= pkg_toStdLogic(false);
      dbus_axi_decoder_io_sharedOutputs_1_arw_rValid <= pkg_toStdLogic(false);
      dbus_axi_decoder_io_input_r_rValid <= pkg_toStdLogic(false);
      axi_ram_io_axi_arbiter_io_output_arw_rValid <= pkg_toStdLogic(false);
      axi_ram_io_axi_arbiter_io_output_w_rValid <= pkg_toStdLogic(false);
      axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rValid <= pkg_toStdLogic(false);
      axi_apbBridge_io_axi_arbiter_io_output_arw_rValid <= pkg_toStdLogic(false);
      axi_apbBridge_io_axi_arbiter_io_output_w_rValid <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      if axi_core_cpu_dBus_cmd_ready = '1' then
        axi_core_cpu_dBus_cmd_rValid <= axi_core_cpu_dBus_cmd_valid;
      end if;
      if axi_core_cpu_dBus_cmd_m2sPipe_ready = '1' then
        axi_core_cpu_dBus_cmd_m2sPipe_rValid <= axi_core_cpu_dBus_cmd_m2sPipe_valid;
      end if;
      if axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_valid = '1' then
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid <= pkg_toStdLogic(true);
      end if;
      if axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready = '1' then
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rValid <= pkg_toStdLogic(false);
      end if;
      zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready <= (zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready + zz_axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_s2mPipe_ready_1);
      if streamFork_3_io_outputs_0_fire = '1' then
        zz_1 <= (not streamFork_3_io_outputs_0_payload_last);
      end if;
      if axi4ReadOnlyDecoder_1_io_outputs_0_ar_valid = '1' then
        axi4ReadOnlyDecoder_1_io_outputs_0_ar_rValid <= pkg_toStdLogic(true);
      end if;
      if axi4ReadOnlyDecoder_1_io_outputs_0_ar_validPipe_fire = '1' then
        axi4ReadOnlyDecoder_1_io_outputs_0_ar_rValid <= pkg_toStdLogic(false);
      end if;
      if dbus_axi_decoder_io_sharedOutputs_0_arw_valid = '1' then
        dbus_axi_decoder_io_sharedOutputs_0_arw_rValid <= pkg_toStdLogic(true);
      end if;
      if dbus_axi_decoder_io_sharedOutputs_0_arw_validPipe_fire = '1' then
        dbus_axi_decoder_io_sharedOutputs_0_arw_rValid <= pkg_toStdLogic(false);
      end if;
      if dbus_axi_decoder_io_sharedOutputs_1_arw_valid = '1' then
        dbus_axi_decoder_io_sharedOutputs_1_arw_rValid <= pkg_toStdLogic(true);
      end if;
      if dbus_axi_decoder_io_sharedOutputs_1_arw_validPipe_fire = '1' then
        dbus_axi_decoder_io_sharedOutputs_1_arw_rValid <= pkg_toStdLogic(false);
      end if;
      if dbus_axi_decoder_io_input_r_ready = '1' then
        dbus_axi_decoder_io_input_r_rValid <= dbus_axi_decoder_io_input_r_valid;
      end if;
      if axi_ram_io_axi_arbiter_io_output_arw_valid = '1' then
        axi_ram_io_axi_arbiter_io_output_arw_rValid <= pkg_toStdLogic(true);
      end if;
      if axi_ram_io_axi_arbiter_io_output_arw_halfPipe_fire = '1' then
        axi_ram_io_axi_arbiter_io_output_arw_rValid <= pkg_toStdLogic(false);
      end if;
      if axi_ram_io_axi_arbiter_io_output_w_valid = '1' then
        axi_ram_io_axi_arbiter_io_output_w_rValid <= pkg_toStdLogic(true);
      end if;
      if axi_ram_io_axi_arbiter_io_output_w_s2mPipe_ready = '1' then
        axi_ram_io_axi_arbiter_io_output_w_rValid <= pkg_toStdLogic(false);
      end if;
      if axi_ram_io_axi_arbiter_io_output_w_s2mPipe_ready = '1' then
        axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rValid <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_valid;
      end if;
      if axi_apbBridge_io_axi_arbiter_io_output_arw_valid = '1' then
        axi_apbBridge_io_axi_arbiter_io_output_arw_rValid <= pkg_toStdLogic(true);
      end if;
      if axi_apbBridge_io_axi_arbiter_io_output_arw_halfPipe_fire = '1' then
        axi_apbBridge_io_axi_arbiter_io_output_arw_rValid <= pkg_toStdLogic(false);
      end if;
      if axi_apbBridge_io_axi_arbiter_io_output_w_valid = '1' then
        axi_apbBridge_io_axi_arbiter_io_output_w_rValid <= pkg_toStdLogic(true);
      end if;
      if axi_apbBridge_io_axi_arbiter_io_output_w_halfPipe_fire = '1' then
        axi_apbBridge_io_axi_arbiter_io_output_w_rValid <= pkg_toStdLogic(false);
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      if axi_core_cpu_dBus_cmd_ready = '1' then
        axi_core_cpu_dBus_cmd_rData_wr <= axi_core_cpu_dBus_cmd_payload_wr;
        axi_core_cpu_dBus_cmd_rData_uncached <= axi_core_cpu_dBus_cmd_payload_uncached;
        axi_core_cpu_dBus_cmd_rData_address <= axi_core_cpu_dBus_cmd_payload_address;
        axi_core_cpu_dBus_cmd_rData_data <= axi_core_cpu_dBus_cmd_payload_data;
        axi_core_cpu_dBus_cmd_rData_mask <= axi_core_cpu_dBus_cmd_payload_mask;
        axi_core_cpu_dBus_cmd_rData_size <= axi_core_cpu_dBus_cmd_payload_size;
        axi_core_cpu_dBus_cmd_rData_last <= axi_core_cpu_dBus_cmd_payload_last;
      end if;
      if axi_core_cpu_dBus_cmd_m2sPipe_ready = '1' then
        axi_core_cpu_dBus_cmd_m2sPipe_rData_wr <= axi_core_cpu_dBus_cmd_m2sPipe_payload_wr;
        axi_core_cpu_dBus_cmd_m2sPipe_rData_uncached <= axi_core_cpu_dBus_cmd_m2sPipe_payload_uncached;
        axi_core_cpu_dBus_cmd_m2sPipe_rData_address <= axi_core_cpu_dBus_cmd_m2sPipe_payload_address;
        axi_core_cpu_dBus_cmd_m2sPipe_rData_data <= axi_core_cpu_dBus_cmd_m2sPipe_payload_data;
        axi_core_cpu_dBus_cmd_m2sPipe_rData_mask <= axi_core_cpu_dBus_cmd_m2sPipe_payload_mask;
        axi_core_cpu_dBus_cmd_m2sPipe_rData_size <= axi_core_cpu_dBus_cmd_m2sPipe_payload_size;
        axi_core_cpu_dBus_cmd_m2sPipe_rData_last <= axi_core_cpu_dBus_cmd_m2sPipe_payload_last;
      end if;
      if axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_ready = '1' then
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_wr <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_wr;
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_uncached <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_uncached;
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_address <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_address;
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_data <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_data;
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_mask <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_mask;
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_size <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_size;
        axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_rData_last <= axi_core_cpu_dBus_cmd_m2sPipe_m2sPipe_payload_last;
      end if;
      if dbus_axi_decoder_io_input_r_ready = '1' then
        dbus_axi_decoder_io_input_r_rData_data <= dbus_axi_decoder_io_input_r_payload_data;
        dbus_axi_decoder_io_input_r_rData_resp <= dbus_axi_decoder_io_input_r_payload_resp;
        dbus_axi_decoder_io_input_r_rData_last <= dbus_axi_decoder_io_input_r_payload_last;
      end if;
      if axi_ram_io_axi_arbiter_io_output_arw_ready = '1' then
        axi_ram_io_axi_arbiter_io_output_arw_rData_addr <= axi_ram_io_axi_arbiter_io_output_arw_payload_addr;
        axi_ram_io_axi_arbiter_io_output_arw_rData_id <= axi_ram_io_axi_arbiter_io_output_arw_payload_id;
        axi_ram_io_axi_arbiter_io_output_arw_rData_len <= axi_ram_io_axi_arbiter_io_output_arw_payload_len;
        axi_ram_io_axi_arbiter_io_output_arw_rData_size <= axi_ram_io_axi_arbiter_io_output_arw_payload_size;
        axi_ram_io_axi_arbiter_io_output_arw_rData_burst <= axi_ram_io_axi_arbiter_io_output_arw_payload_burst;
        axi_ram_io_axi_arbiter_io_output_arw_rData_write <= axi_ram_io_axi_arbiter_io_output_arw_payload_write;
      end if;
      if axi_ram_io_axi_arbiter_io_output_w_ready = '1' then
        axi_ram_io_axi_arbiter_io_output_w_rData_data <= axi_ram_io_axi_arbiter_io_output_w_payload_data;
        axi_ram_io_axi_arbiter_io_output_w_rData_strb <= axi_ram_io_axi_arbiter_io_output_w_payload_strb;
        axi_ram_io_axi_arbiter_io_output_w_rData_last <= axi_ram_io_axi_arbiter_io_output_w_payload_last;
      end if;
      if axi_ram_io_axi_arbiter_io_output_w_s2mPipe_ready = '1' then
        axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_data <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_data;
        axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_strb <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_strb;
        axi_ram_io_axi_arbiter_io_output_w_s2mPipe_rData_last <= axi_ram_io_axi_arbiter_io_output_w_s2mPipe_payload_last;
      end if;
      if axi_apbBridge_io_axi_arbiter_io_output_arw_ready = '1' then
        axi_apbBridge_io_axi_arbiter_io_output_arw_rData_addr <= axi_apbBridge_io_axi_arbiter_io_output_arw_payload_addr;
        axi_apbBridge_io_axi_arbiter_io_output_arw_rData_id <= axi_apbBridge_io_axi_arbiter_io_output_arw_payload_id;
        axi_apbBridge_io_axi_arbiter_io_output_arw_rData_len <= axi_apbBridge_io_axi_arbiter_io_output_arw_payload_len;
        axi_apbBridge_io_axi_arbiter_io_output_arw_rData_size <= axi_apbBridge_io_axi_arbiter_io_output_arw_payload_size;
        axi_apbBridge_io_axi_arbiter_io_output_arw_rData_burst <= axi_apbBridge_io_axi_arbiter_io_output_arw_payload_burst;
        axi_apbBridge_io_axi_arbiter_io_output_arw_rData_write <= axi_apbBridge_io_axi_arbiter_io_output_arw_payload_write;
      end if;
      if axi_apbBridge_io_axi_arbiter_io_output_w_ready = '1' then
        axi_apbBridge_io_axi_arbiter_io_output_w_rData_data <= axi_apbBridge_io_axi_arbiter_io_output_w_payload_data;
        axi_apbBridge_io_axi_arbiter_io_output_w_rData_strb <= axi_apbBridge_io_axi_arbiter_io_output_w_payload_strb;
        axi_apbBridge_io_axi_arbiter_io_output_w_rData_last <= axi_apbBridge_io_axi_arbiter_io_output_w_payload_last;
      end if;
    end if;
  end process;

  process(io_mainClk)
  begin
    if rising_edge(io_mainClk) then
      axi_core_cpu_debug_resetOut_regNext <= axi_core_cpu_debug_resetOut;
    end if;
  end process;

  process(io_mainClk, resetCtrl_systemReset)
  begin
    if resetCtrl_systemReset = '1' then
      axi_core_cpu_debug_bus_cmd_fire_regNext <= pkg_toStdLogic(false);
    elsif rising_edge(io_mainClk) then
      axi_core_cpu_debug_bus_cmd_fire_regNext <= axi_core_cpu_debug_bus_cmd_fire;
    end if;
  end process;

end arch;

